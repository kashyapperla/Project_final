
module fpalu_add1_DW01_inc_0 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[7]), .IN2(A[7]), .Q(SUM[7]) );
endmodule


module fpalu_add1_DW01_sub_22 ( A, B, CI, DIFF, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  NOR2X0 U1 ( .IN1(B[1]), .IN2(\B[0] ), .QN(n21) );
  AND2X1 U2 ( .IN1(n44), .IN2(n21), .Q(n1) );
  AND2X1 U3 ( .IN1(n43), .IN2(n1), .Q(n2) );
  AND2X1 U4 ( .IN1(n42), .IN2(n2), .Q(n3) );
  AND2X1 U5 ( .IN1(n41), .IN2(n3), .Q(n4) );
  AND2X1 U6 ( .IN1(n40), .IN2(n4), .Q(n5) );
  AND2X1 U7 ( .IN1(n39), .IN2(n5), .Q(n6) );
  AND2X1 U8 ( .IN1(n38), .IN2(n6), .Q(n7) );
  AND2X1 U9 ( .IN1(n37), .IN2(n7), .Q(n8) );
  AND2X1 U10 ( .IN1(n36), .IN2(n8), .Q(n9) );
  AND2X1 U11 ( .IN1(n35), .IN2(n9), .Q(n10) );
  AND2X1 U12 ( .IN1(n34), .IN2(n10), .Q(n11) );
  AND2X1 U13 ( .IN1(n33), .IN2(n11), .Q(n12) );
  AND2X1 U14 ( .IN1(n32), .IN2(n12), .Q(n13) );
  AND2X1 U15 ( .IN1(n31), .IN2(n13), .Q(n14) );
  AND2X1 U16 ( .IN1(n30), .IN2(n14), .Q(n15) );
  AND2X1 U17 ( .IN1(n29), .IN2(n15), .Q(n16) );
  AND2X1 U18 ( .IN1(n28), .IN2(n16), .Q(n17) );
  AND2X1 U19 ( .IN1(n27), .IN2(n17), .Q(n18) );
  AND2X1 U20 ( .IN1(n26), .IN2(n18), .Q(n19) );
  AND2X1 U21 ( .IN1(n25), .IN2(n19), .Q(n20) );
  NAND2X1 U22 ( .IN1(n24), .IN2(n20), .QN(n22) );
  INVX0 U23 ( .INP(B[1]), .ZN(n45) );
  INVX0 U24 ( .INP(B[2]), .ZN(n44) );
  INVX0 U25 ( .INP(B[3]), .ZN(n43) );
  INVX0 U26 ( .INP(B[4]), .ZN(n42) );
  INVX0 U27 ( .INP(B[5]), .ZN(n41) );
  INVX0 U28 ( .INP(B[6]), .ZN(n40) );
  INVX0 U29 ( .INP(B[7]), .ZN(n39) );
  INVX0 U30 ( .INP(B[8]), .ZN(n38) );
  INVX0 U31 ( .INP(B[9]), .ZN(n37) );
  INVX0 U32 ( .INP(B[10]), .ZN(n36) );
  INVX0 U33 ( .INP(B[11]), .ZN(n35) );
  INVX0 U34 ( .INP(B[12]), .ZN(n34) );
  INVX0 U35 ( .INP(B[13]), .ZN(n33) );
  INVX0 U36 ( .INP(B[14]), .ZN(n32) );
  INVX0 U37 ( .INP(B[15]), .ZN(n31) );
  INVX0 U38 ( .INP(B[16]), .ZN(n30) );
  INVX0 U39 ( .INP(B[17]), .ZN(n29) );
  INVX0 U40 ( .INP(B[18]), .ZN(n28) );
  INVX0 U41 ( .INP(B[19]), .ZN(n27) );
  INVX0 U42 ( .INP(B[20]), .ZN(n26) );
  INVX0 U43 ( .INP(B[21]), .ZN(n25) );
  INVX0 U44 ( .INP(B[22]), .ZN(n24) );
  INVX0 U45 ( .INP(\B[0] ), .ZN(n46) );
  XNOR2X1 U46 ( .IN1(n23), .IN2(n22), .Q(DIFF[23]) );
  INVX0 U47 ( .INP(B[23]), .ZN(n23) );
  XOR2X1 U48 ( .IN1(n24), .IN2(n20), .Q(DIFF[22]) );
  XOR2X1 U49 ( .IN1(n25), .IN2(n19), .Q(DIFF[21]) );
  XOR2X1 U50 ( .IN1(n26), .IN2(n18), .Q(DIFF[20]) );
  XOR2X1 U51 ( .IN1(n27), .IN2(n17), .Q(DIFF[19]) );
  XOR2X1 U52 ( .IN1(n28), .IN2(n16), .Q(DIFF[18]) );
  XOR2X1 U53 ( .IN1(n29), .IN2(n15), .Q(DIFF[17]) );
  XOR2X1 U54 ( .IN1(n30), .IN2(n14), .Q(DIFF[16]) );
  XOR2X1 U55 ( .IN1(n31), .IN2(n13), .Q(DIFF[15]) );
  XOR2X1 U56 ( .IN1(n32), .IN2(n12), .Q(DIFF[14]) );
  XOR2X1 U57 ( .IN1(n33), .IN2(n11), .Q(DIFF[13]) );
  XOR2X1 U58 ( .IN1(n34), .IN2(n10), .Q(DIFF[12]) );
  XOR2X1 U59 ( .IN1(n35), .IN2(n9), .Q(DIFF[11]) );
  XOR2X1 U60 ( .IN1(n36), .IN2(n8), .Q(DIFF[10]) );
  XOR2X1 U61 ( .IN1(n37), .IN2(n7), .Q(DIFF[9]) );
  XOR2X1 U62 ( .IN1(n38), .IN2(n6), .Q(DIFF[8]) );
  XOR2X1 U63 ( .IN1(n39), .IN2(n5), .Q(DIFF[7]) );
  XOR2X1 U64 ( .IN1(n40), .IN2(n4), .Q(DIFF[6]) );
  XOR2X1 U65 ( .IN1(n41), .IN2(n3), .Q(DIFF[5]) );
  XOR2X1 U66 ( .IN1(n42), .IN2(n2), .Q(DIFF[4]) );
  XOR2X1 U67 ( .IN1(n43), .IN2(n1), .Q(DIFF[3]) );
  XOR2X1 U68 ( .IN1(n44), .IN2(n21), .Q(DIFF[2]) );
  XOR2X1 U69 ( .IN1(n45), .IN2(n46), .Q(DIFF[1]) );
endmodule


module fpalu_add1_DW01_add_0 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [23:1] carry;

  FADDX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FADDX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  FADDX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  FADDX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FADDX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  FADDX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X1 U1_23 ( .IN1(A[23]), .IN2(B[23]), .IN3(carry[23]), .Q(SUM[23]) );
  AND2X1 U1 ( .IN1(A[0]), .IN2(B[0]), .Q(n1) );
  XOR2X1 U2 ( .IN1(A[0]), .IN2(B[0]), .Q(SUM[0]) );
endmodule


module fpalu_add1_DW01_add_1 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [23:1] carry;

  FADDX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FADDX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  FADDX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  FADDX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FADDX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  FADDX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  INVX0 U1 ( .INP(carry[23]), .ZN(n2) );
  AND2X1 U2 ( .IN1(A[0]), .IN2(B[0]), .Q(n1) );
  XOR2X1 U3 ( .IN1(n2), .IN2(B[23]), .Q(SUM[23]) );
  XOR2X1 U4 ( .IN1(A[0]), .IN2(B[0]), .Q(SUM[0]) );
endmodule


module fpalu_add1_DW01_sub_23 ( A, B, CI, DIFF, CO );
  input [24:0] A;
  input [24:0] B;
  output [24:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  NOR2X0 U1 ( .IN1(B[1]), .IN2(\B[0] ), .QN(n21) );
  AND2X1 U2 ( .IN1(n41), .IN2(n4), .Q(n1) );
  AND2X1 U3 ( .IN1(n39), .IN2(n10), .Q(n2) );
  AND2X1 U4 ( .IN1(n42), .IN2(n1), .Q(n3) );
  AND2X1 U5 ( .IN1(n40), .IN2(n2), .Q(n4) );
  INVX0 U6 ( .INP(B[22]), .ZN(n43) );
  INVX0 U7 ( .INP(B[16]), .ZN(n39) );
  INVX0 U8 ( .INP(B[17]), .ZN(n40) );
  INVX0 U9 ( .INP(B[18]), .ZN(n41) );
  INVX0 U10 ( .INP(B[19]), .ZN(n42) );
  AND2X1 U11 ( .IN1(n37), .IN2(n16), .Q(n5) );
  AND2X1 U12 ( .IN1(n31), .IN2(n14), .Q(n6) );
  AND2X1 U13 ( .IN1(n38), .IN2(n5), .Q(n7) );
  AND2X1 U14 ( .IN1(n32), .IN2(n6), .Q(n8) );
  AND2X1 U15 ( .IN1(n33), .IN2(n8), .Q(n9) );
  AND2X1 U16 ( .IN1(n34), .IN2(n9), .Q(n10) );
  AND2X1 U17 ( .IN1(n29), .IN2(n7), .Q(n11) );
  AND2X1 U18 ( .IN1(n23), .IN2(n20), .Q(n12) );
  AND2X1 U19 ( .IN1(n26), .IN2(n15), .Q(n13) );
  AND2X1 U20 ( .IN1(n30), .IN2(n11), .Q(n14) );
  AND2X1 U21 ( .IN1(n24), .IN2(n12), .Q(n15) );
  AND2X1 U22 ( .IN1(n25), .IN2(n13), .Q(n16) );
  AND2X1 U23 ( .IN1(n35), .IN2(n3), .Q(n17) );
  AND2X1 U24 ( .IN1(n36), .IN2(n17), .Q(n18) );
  INVX0 U25 ( .INP(B[8]), .ZN(n37) );
  INVX0 U26 ( .INP(B[12]), .ZN(n31) );
  INVX0 U27 ( .INP(B[9]), .ZN(n38) );
  INVX0 U28 ( .INP(B[13]), .ZN(n32) );
  INVX0 U29 ( .INP(B[15]), .ZN(n34) );
  INVX0 U30 ( .INP(B[14]), .ZN(n33) );
  INVX0 U31 ( .INP(B[10]), .ZN(n29) );
  INVX0 U32 ( .INP(B[4]), .ZN(n23) );
  INVX0 U33 ( .INP(B[6]), .ZN(n26) );
  INVX0 U34 ( .INP(B[11]), .ZN(n30) );
  INVX0 U35 ( .INP(B[5]), .ZN(n24) );
  INVX0 U36 ( .INP(B[7]), .ZN(n25) );
  INVX0 U37 ( .INP(B[20]), .ZN(n35) );
  INVX0 U38 ( .INP(B[1]), .ZN(n44) );
  INVX0 U39 ( .INP(B[21]), .ZN(n36) );
  AND2X1 U40 ( .IN1(n28), .IN2(n21), .Q(n19) );
  AND2X1 U41 ( .IN1(n27), .IN2(n19), .Q(n20) );
  XOR2X1 U42 ( .IN1(B[23]), .IN2(n22), .Q(DIFF[23]) );
  NAND2X1 U43 ( .IN1(n43), .IN2(n18), .QN(n22) );
  INVX0 U44 ( .INP(B[2]), .ZN(n28) );
  INVX0 U45 ( .INP(B[3]), .ZN(n27) );
  INVX0 U46 ( .INP(\B[0] ), .ZN(n45) );
  XOR2X1 U47 ( .IN1(n43), .IN2(n18), .Q(DIFF[22]) );
  XOR2X1 U48 ( .IN1(n36), .IN2(n17), .Q(DIFF[21]) );
  XOR2X1 U49 ( .IN1(n35), .IN2(n3), .Q(DIFF[20]) );
  XOR2X1 U50 ( .IN1(n42), .IN2(n1), .Q(DIFF[19]) );
  XOR2X1 U51 ( .IN1(n41), .IN2(n4), .Q(DIFF[18]) );
  XOR2X1 U52 ( .IN1(n40), .IN2(n2), .Q(DIFF[17]) );
  XOR2X1 U53 ( .IN1(n39), .IN2(n10), .Q(DIFF[16]) );
  XOR2X1 U54 ( .IN1(n34), .IN2(n9), .Q(DIFF[15]) );
  XOR2X1 U55 ( .IN1(n33), .IN2(n8), .Q(DIFF[14]) );
  XOR2X1 U56 ( .IN1(n32), .IN2(n6), .Q(DIFF[13]) );
  XOR2X1 U57 ( .IN1(n31), .IN2(n14), .Q(DIFF[12]) );
  XOR2X1 U58 ( .IN1(n30), .IN2(n11), .Q(DIFF[11]) );
  XOR2X1 U59 ( .IN1(n29), .IN2(n7), .Q(DIFF[10]) );
  XOR2X1 U60 ( .IN1(n38), .IN2(n5), .Q(DIFF[9]) );
  XOR2X1 U61 ( .IN1(n37), .IN2(n16), .Q(DIFF[8]) );
  XOR2X1 U62 ( .IN1(n25), .IN2(n13), .Q(DIFF[7]) );
  XOR2X1 U63 ( .IN1(n26), .IN2(n15), .Q(DIFF[6]) );
  XOR2X1 U64 ( .IN1(n24), .IN2(n12), .Q(DIFF[5]) );
  XOR2X1 U65 ( .IN1(n23), .IN2(n20), .Q(DIFF[4]) );
  XOR2X1 U66 ( .IN1(n27), .IN2(n19), .Q(DIFF[3]) );
  XOR2X1 U67 ( .IN1(n28), .IN2(n21), .Q(DIFF[2]) );
  XOR2X1 U68 ( .IN1(n44), .IN2(n45), .Q(DIFF[1]) );
endmodule


module fpalu_add1_DW01_sub_24 ( A, B, CI, DIFF, CO );
  input [24:0] A;
  input [24:0] B;
  output [24:0] DIFF;
  input CI;
  output CO;
  wire   \B[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45;
  assign DIFF[0] = \B[0] ;
  assign \B[0]  = B[0];

  NOR2X0 U1 ( .IN1(B[1]), .IN2(\B[0] ), .QN(n1) );
  AND2X1 U2 ( .IN1(n39), .IN2(n12), .Q(n2) );
  AND2X1 U3 ( .IN1(n41), .IN2(n13), .Q(n3) );
  AND2X1 U4 ( .IN1(n43), .IN2(n14), .Q(n4) );
  AND2X1 U5 ( .IN1(n45), .IN2(n15), .Q(n5) );
  AND2X1 U6 ( .IN1(n25), .IN2(n16), .Q(n6) );
  AND2X1 U7 ( .IN1(n27), .IN2(n17), .Q(n7) );
  AND2X1 U8 ( .IN1(n29), .IN2(n18), .Q(n8) );
  AND2X1 U9 ( .IN1(n31), .IN2(n19), .Q(n9) );
  AND2X1 U10 ( .IN1(n33), .IN2(n20), .Q(n10) );
  AND2X1 U11 ( .IN1(n36), .IN2(n21), .Q(n11) );
  AND2X1 U12 ( .IN1(n38), .IN2(n1), .Q(n12) );
  AND2X1 U13 ( .IN1(n40), .IN2(n2), .Q(n13) );
  AND2X1 U14 ( .IN1(n42), .IN2(n3), .Q(n14) );
  AND2X1 U15 ( .IN1(n44), .IN2(n4), .Q(n15) );
  AND2X1 U16 ( .IN1(n24), .IN2(n5), .Q(n16) );
  AND2X1 U17 ( .IN1(n26), .IN2(n6), .Q(n17) );
  AND2X1 U18 ( .IN1(n28), .IN2(n7), .Q(n18) );
  AND2X1 U19 ( .IN1(n30), .IN2(n8), .Q(n19) );
  AND2X1 U20 ( .IN1(n32), .IN2(n9), .Q(n20) );
  AND2X1 U21 ( .IN1(n35), .IN2(n10), .Q(n21) );
  AND2X1 U22 ( .IN1(n37), .IN2(n11), .Q(DIFF[23]) );
  INVX0 U23 ( .INP(B[22]), .ZN(n37) );
  INVX0 U24 ( .INP(B[1]), .ZN(n34) );
  INVX0 U25 ( .INP(B[3]), .ZN(n39) );
  INVX0 U26 ( .INP(B[5]), .ZN(n41) );
  INVX0 U27 ( .INP(B[7]), .ZN(n43) );
  INVX0 U28 ( .INP(B[9]), .ZN(n45) );
  INVX0 U29 ( .INP(B[11]), .ZN(n25) );
  INVX0 U30 ( .INP(B[13]), .ZN(n27) );
  INVX0 U31 ( .INP(B[15]), .ZN(n29) );
  INVX0 U32 ( .INP(B[17]), .ZN(n31) );
  INVX0 U33 ( .INP(B[19]), .ZN(n33) );
  INVX0 U34 ( .INP(B[21]), .ZN(n36) );
  INVX0 U35 ( .INP(B[2]), .ZN(n38) );
  INVX0 U36 ( .INP(B[4]), .ZN(n40) );
  INVX0 U37 ( .INP(B[6]), .ZN(n42) );
  INVX0 U38 ( .INP(B[8]), .ZN(n44) );
  INVX0 U39 ( .INP(B[10]), .ZN(n24) );
  INVX0 U40 ( .INP(B[12]), .ZN(n26) );
  INVX0 U41 ( .INP(B[14]), .ZN(n28) );
  INVX0 U42 ( .INP(B[16]), .ZN(n30) );
  INVX0 U43 ( .INP(B[18]), .ZN(n32) );
  INVX0 U44 ( .INP(B[20]), .ZN(n35) );
  INVX0 U45 ( .INP(\B[0] ), .ZN(n23) );
  XOR2X1 U46 ( .IN1(n37), .IN2(n11), .Q(DIFF[22]) );
  XOR2X1 U47 ( .IN1(n36), .IN2(n21), .Q(DIFF[21]) );
  XOR2X1 U48 ( .IN1(n35), .IN2(n10), .Q(DIFF[20]) );
  XOR2X1 U49 ( .IN1(n33), .IN2(n20), .Q(DIFF[19]) );
  XOR2X1 U50 ( .IN1(n32), .IN2(n9), .Q(DIFF[18]) );
  XOR2X1 U51 ( .IN1(n31), .IN2(n19), .Q(DIFF[17]) );
  XOR2X1 U52 ( .IN1(n30), .IN2(n8), .Q(DIFF[16]) );
  XOR2X1 U53 ( .IN1(n29), .IN2(n18), .Q(DIFF[15]) );
  XOR2X1 U54 ( .IN1(n28), .IN2(n7), .Q(DIFF[14]) );
  XOR2X1 U55 ( .IN1(n27), .IN2(n17), .Q(DIFF[13]) );
  XOR2X1 U56 ( .IN1(n26), .IN2(n6), .Q(DIFF[12]) );
  XOR2X1 U57 ( .IN1(n25), .IN2(n16), .Q(DIFF[11]) );
  XOR2X1 U58 ( .IN1(n24), .IN2(n5), .Q(DIFF[10]) );
  XOR2X1 U59 ( .IN1(n45), .IN2(n15), .Q(DIFF[9]) );
  XOR2X1 U60 ( .IN1(n44), .IN2(n4), .Q(DIFF[8]) );
  XOR2X1 U61 ( .IN1(n43), .IN2(n14), .Q(DIFF[7]) );
  XOR2X1 U62 ( .IN1(n42), .IN2(n3), .Q(DIFF[6]) );
  XOR2X1 U63 ( .IN1(n41), .IN2(n13), .Q(DIFF[5]) );
  XOR2X1 U64 ( .IN1(n40), .IN2(n2), .Q(DIFF[4]) );
  XOR2X1 U65 ( .IN1(n39), .IN2(n12), .Q(DIFF[3]) );
  XOR2X1 U66 ( .IN1(n38), .IN2(n1), .Q(DIFF[2]) );
  XOR2X1 U67 ( .IN1(n34), .IN2(n23), .Q(DIFF[1]) );
endmodule


module fpalu_add1_DW01_add_2 ( A, B, CI, SUM, CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [23:1] carry;

  FADDX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FADDX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  FADDX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  FADDX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FADDX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  FADDX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  INVX0 U1 ( .INP(carry[23]), .ZN(n2) );
  AND2X1 U2 ( .IN1(A[0]), .IN2(B[0]), .Q(n1) );
  XOR2X1 U3 ( .IN1(n2), .IN2(B[23]), .Q(SUM[23]) );
  XOR2X1 U4 ( .IN1(A[0]), .IN2(B[0]), .Q(SUM[0]) );
endmodule


module fpalu_add1_DW01_cmp6_0 ( A, B, TC, LT, GT, EQ, LE, GE, NE );
  input [25:0] A;
  input [25:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125;

  INVX0 U1 ( .INP(B[22]), .ZN(n13) );
  INVX0 U2 ( .INP(B[17]), .ZN(n11) );
  INVX0 U3 ( .INP(B[19]), .ZN(n12) );
  INVX0 U4 ( .INP(B[9]), .ZN(n10) );
  INVX0 U5 ( .INP(B[13]), .ZN(n5) );
  INVX0 U6 ( .INP(B[15]), .ZN(n6) );
  INVX0 U7 ( .INP(B[11]), .ZN(n4) );
  INVX0 U8 ( .INP(B[5]), .ZN(n1) );
  INVX0 U9 ( .INP(B[7]), .ZN(n2) );
  INVX0 U10 ( .INP(B[21]), .ZN(n8) );
  INVX0 U11 ( .INP(B[23]), .ZN(n9) );
  INVX0 U12 ( .INP(B[1]), .ZN(n14) );
  INVX0 U13 ( .INP(B[3]), .ZN(n3) );
  INVX0 U14 ( .INP(B[0]), .ZN(n16) );
  INVX0 U15 ( .INP(n92), .ZN(n15) );
  INVX0 U16 ( .INP(A[1]), .ZN(n22) );
  INVX0 U17 ( .INP(A[2]), .ZN(n24) );
  INVX0 U18 ( .INP(A[4]), .ZN(n25) );
  INVX0 U19 ( .INP(A[6]), .ZN(n26) );
  INVX0 U20 ( .INP(A[8]), .ZN(n27) );
  INVX0 U21 ( .INP(A[10]), .ZN(n17) );
  INVX0 U22 ( .INP(A[12]), .ZN(n18) );
  INVX0 U23 ( .INP(A[14]), .ZN(n19) );
  INVX0 U24 ( .INP(A[16]), .ZN(n20) );
  INVX0 U25 ( .INP(A[18]), .ZN(n21) );
  INVX0 U26 ( .INP(A[20]), .ZN(n23) );
  INVX0 U27 ( .INP(n35), .ZN(n7) );
  NOR2X0 U28 ( .IN1(n28), .IN2(n9), .QN(LT) );
  OA21X1 U29 ( .IN1(A[22]), .IN2(n13), .IN3(n29), .Q(n28) );
  NAND3X0 U30 ( .IN1(n30), .IN2(n31), .IN3(n32), .QN(n29) );
  NAND3X0 U31 ( .IN1(n33), .IN2(n34), .IN3(n7), .QN(n30) );
  NAND3X0 U32 ( .IN1(n36), .IN2(n37), .IN3(n38), .QN(n33) );
  NAND3X0 U33 ( .IN1(n39), .IN2(n40), .IN3(n41), .QN(n36) );
  NAND3X0 U34 ( .IN1(n42), .IN2(n43), .IN3(n44), .QN(n39) );
  NAND3X0 U35 ( .IN1(n45), .IN2(n46), .IN3(n47), .QN(n42) );
  NAND3X0 U36 ( .IN1(n48), .IN2(n49), .IN3(n50), .QN(n45) );
  NAND3X0 U37 ( .IN1(n51), .IN2(n52), .IN3(n53), .QN(n48) );
  NAND3X0 U38 ( .IN1(n54), .IN2(n55), .IN3(n56), .QN(n51) );
  NAND3X0 U39 ( .IN1(n57), .IN2(n58), .IN3(n59), .QN(n54) );
  NAND3X0 U40 ( .IN1(n60), .IN2(n61), .IN3(n62), .QN(n57) );
  NAND3X0 U41 ( .IN1(n63), .IN2(n64), .IN3(n65), .QN(n60) );
  NAND3X0 U42 ( .IN1(n66), .IN2(n67), .IN3(n68), .QN(n63) );
  NAND3X0 U43 ( .IN1(n69), .IN2(n70), .IN3(n71), .QN(n66) );
  NAND3X0 U44 ( .IN1(n72), .IN2(n73), .IN3(n74), .QN(n69) );
  NAND3X0 U45 ( .IN1(n75), .IN2(n76), .IN3(n77), .QN(n72) );
  NAND3X0 U46 ( .IN1(n78), .IN2(n79), .IN3(n80), .QN(n75) );
  NAND3X0 U47 ( .IN1(n81), .IN2(n82), .IN3(n83), .QN(n78) );
  NAND3X0 U48 ( .IN1(n84), .IN2(n85), .IN3(n86), .QN(n81) );
  NAND3X0 U49 ( .IN1(n87), .IN2(n88), .IN3(n89), .QN(n84) );
  AO221X1 U50 ( .IN1(n90), .IN2(n14), .IN3(A[1]), .IN4(n15), .IN5(n91), .Q(n87) );
  NAND2X0 U51 ( .IN1(n92), .IN2(n22), .QN(n90) );
  NOR2X0 U52 ( .IN1(n16), .IN2(A[0]), .QN(n92) );
  AO221X1 U53 ( .IN1(n93), .IN2(n32), .IN3(A[22]), .IN4(n13), .IN5(n9), .Q(GT)
         );
  XNOR2X1 U54 ( .IN1(A[22]), .IN2(B[22]), .Q(n32) );
  NOR2X0 U55 ( .IN1(n35), .IN2(n94), .QN(n93) );
  AND3X1 U56 ( .IN1(n31), .IN2(n95), .IN3(n96), .Q(n94) );
  NAND3X0 U57 ( .IN1(n97), .IN2(n41), .IN3(n38), .QN(n96) );
  AND2X1 U58 ( .IN1(n95), .IN2(n34), .Q(n38) );
  NAND2X0 U59 ( .IN1(B[20]), .IN2(n23), .QN(n34) );
  OR2X1 U60 ( .IN1(n12), .IN2(A[19]), .Q(n41) );
  NAND3X0 U61 ( .IN1(n37), .IN2(n98), .IN3(n99), .QN(n97) );
  NAND3X0 U62 ( .IN1(n100), .IN2(n47), .IN3(n44), .QN(n99) );
  AND2X1 U63 ( .IN1(n98), .IN2(n40), .Q(n44) );
  NAND2X0 U64 ( .IN1(B[18]), .IN2(n21), .QN(n40) );
  OR2X1 U65 ( .IN1(n11), .IN2(A[17]), .Q(n47) );
  NAND3X0 U66 ( .IN1(n43), .IN2(n101), .IN3(n102), .QN(n100) );
  NAND3X0 U67 ( .IN1(n103), .IN2(n53), .IN3(n50), .QN(n102) );
  AND2X1 U68 ( .IN1(n101), .IN2(n46), .Q(n50) );
  NAND2X0 U69 ( .IN1(B[16]), .IN2(n20), .QN(n46) );
  OR2X1 U70 ( .IN1(n6), .IN2(A[15]), .Q(n53) );
  NAND3X0 U71 ( .IN1(n49), .IN2(n104), .IN3(n105), .QN(n103) );
  NAND3X0 U72 ( .IN1(n106), .IN2(n59), .IN3(n56), .QN(n105) );
  AND2X1 U73 ( .IN1(n104), .IN2(n52), .Q(n56) );
  NAND2X0 U74 ( .IN1(B[14]), .IN2(n19), .QN(n52) );
  OR2X1 U75 ( .IN1(n5), .IN2(A[13]), .Q(n59) );
  NAND3X0 U76 ( .IN1(n55), .IN2(n107), .IN3(n108), .QN(n106) );
  NAND3X0 U77 ( .IN1(n109), .IN2(n65), .IN3(n62), .QN(n108) );
  AND2X1 U78 ( .IN1(n107), .IN2(n58), .Q(n62) );
  NAND2X0 U79 ( .IN1(B[12]), .IN2(n18), .QN(n58) );
  OR2X1 U80 ( .IN1(n4), .IN2(A[11]), .Q(n65) );
  NAND3X0 U81 ( .IN1(n61), .IN2(n110), .IN3(n111), .QN(n109) );
  NAND3X0 U82 ( .IN1(n112), .IN2(n71), .IN3(n68), .QN(n111) );
  AND2X1 U83 ( .IN1(n110), .IN2(n64), .Q(n68) );
  NAND2X0 U84 ( .IN1(B[10]), .IN2(n17), .QN(n64) );
  OR2X1 U85 ( .IN1(n10), .IN2(A[9]), .Q(n71) );
  NAND3X0 U86 ( .IN1(n67), .IN2(n113), .IN3(n114), .QN(n112) );
  NAND3X0 U87 ( .IN1(n115), .IN2(n77), .IN3(n74), .QN(n114) );
  AND2X1 U88 ( .IN1(n113), .IN2(n70), .Q(n74) );
  NAND2X0 U89 ( .IN1(B[8]), .IN2(n27), .QN(n70) );
  OR2X1 U90 ( .IN1(n2), .IN2(A[7]), .Q(n77) );
  NAND3X0 U91 ( .IN1(n73), .IN2(n116), .IN3(n117), .QN(n115) );
  NAND3X0 U92 ( .IN1(n118), .IN2(n83), .IN3(n80), .QN(n117) );
  AND2X1 U93 ( .IN1(n116), .IN2(n76), .Q(n80) );
  NAND2X0 U94 ( .IN1(B[6]), .IN2(n26), .QN(n76) );
  OR2X1 U95 ( .IN1(n1), .IN2(A[5]), .Q(n83) );
  NAND3X0 U96 ( .IN1(n79), .IN2(n119), .IN3(n120), .QN(n118) );
  NAND3X0 U97 ( .IN1(n121), .IN2(n89), .IN3(n86), .QN(n120) );
  AND2X1 U98 ( .IN1(n119), .IN2(n82), .Q(n86) );
  NAND2X0 U99 ( .IN1(B[4]), .IN2(n25), .QN(n82) );
  OR2X1 U100 ( .IN1(n3), .IN2(A[3]), .Q(n89) );
  NAND3X0 U101 ( .IN1(n85), .IN2(n122), .IN3(n123), .QN(n121) );
  AO221X1 U102 ( .IN1(B[1]), .IN2(n124), .IN3(n125), .IN4(n22), .IN5(n91), .Q(
        n123) );
  NAND2X0 U103 ( .IN1(n122), .IN2(n88), .QN(n91) );
  NAND2X0 U104 ( .IN1(B[2]), .IN2(n24), .QN(n88) );
  OR2X1 U105 ( .IN1(n125), .IN2(n22), .Q(n124) );
  NAND2X0 U106 ( .IN1(A[0]), .IN2(n16), .QN(n125) );
  OR2X1 U107 ( .IN1(n24), .IN2(B[2]), .Q(n122) );
  NAND2X0 U108 ( .IN1(A[3]), .IN2(n3), .QN(n85) );
  OR2X1 U109 ( .IN1(n25), .IN2(B[4]), .Q(n119) );
  NAND2X0 U110 ( .IN1(A[5]), .IN2(n1), .QN(n79) );
  OR2X1 U111 ( .IN1(n26), .IN2(B[6]), .Q(n116) );
  NAND2X0 U112 ( .IN1(A[7]), .IN2(n2), .QN(n73) );
  OR2X1 U113 ( .IN1(n27), .IN2(B[8]), .Q(n113) );
  NAND2X0 U114 ( .IN1(A[9]), .IN2(n10), .QN(n67) );
  OR2X1 U115 ( .IN1(n17), .IN2(B[10]), .Q(n110) );
  NAND2X0 U116 ( .IN1(A[11]), .IN2(n4), .QN(n61) );
  OR2X1 U117 ( .IN1(n18), .IN2(B[12]), .Q(n107) );
  NAND2X0 U118 ( .IN1(A[13]), .IN2(n5), .QN(n55) );
  OR2X1 U119 ( .IN1(n19), .IN2(B[14]), .Q(n104) );
  NAND2X0 U120 ( .IN1(A[15]), .IN2(n6), .QN(n49) );
  OR2X1 U121 ( .IN1(n20), .IN2(B[16]), .Q(n101) );
  NAND2X0 U122 ( .IN1(A[17]), .IN2(n11), .QN(n43) );
  OR2X1 U123 ( .IN1(n21), .IN2(B[18]), .Q(n98) );
  NAND2X0 U124 ( .IN1(A[19]), .IN2(n12), .QN(n37) );
  OR2X1 U125 ( .IN1(n23), .IN2(B[20]), .Q(n95) );
  NAND2X0 U126 ( .IN1(A[21]), .IN2(n8), .QN(n31) );
  NOR2X0 U127 ( .IN1(n8), .IN2(A[21]), .QN(n35) );
endmodule


module fpalu_add1_DW_rash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [23:0] A;
  input [7:0] SH;
  output [23:0] B;
  input DATA_TC, SH_TC;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104;

  NAND3X0 U3 ( .IN1(n65), .IN2(n66), .IN3(n1), .QN(n69) );
  INVX0 U4 ( .INP(n55), .ZN(n10) );
  INVX0 U5 ( .INP(n79), .ZN(n13) );
  INVX0 U6 ( .INP(n56), .ZN(n9) );
  INVX0 U7 ( .INP(n78), .ZN(n12) );
  INVX0 U8 ( .INP(n68), .ZN(n7) );
  INVX0 U9 ( .INP(n75), .ZN(n4) );
  INVX0 U10 ( .INP(n66), .ZN(n2) );
  INVX0 U11 ( .INP(n91), .ZN(n3) );
  INVX0 U12 ( .INP(SH[0]), .ZN(n14) );
  INVX0 U13 ( .INP(SH[1]), .ZN(n11) );
  INVX0 U14 ( .INP(n80), .ZN(n5) );
  INVX0 U15 ( .INP(n82), .ZN(n6) );
  NOR2X0 U16 ( .IN1(SH[3]), .IN2(n103), .QN(n65) );
  INVX0 U17 ( .INP(SH[2]), .ZN(n8) );
  INVX0 U18 ( .INP(A[1]), .ZN(n15) );
  INVX0 U19 ( .INP(SH[7]), .ZN(n1) );
  INVX0 U20 ( .INP(A[4]), .ZN(n18) );
  INVX0 U21 ( .INP(A[3]), .ZN(n17) );
  INVX0 U22 ( .INP(A[2]), .ZN(n16) );
  AO222X1 U23 ( .IN1(n19), .IN2(n20), .IN3(n21), .IN4(n22), .IN5(n23), .IN6(
        n24), .Q(B[9]) );
  AO222X1 U24 ( .IN1(n19), .IN2(n25), .IN3(n21), .IN4(n26), .IN5(n23), .IN6(
        n27), .Q(B[8]) );
  AO221X1 U25 ( .IN1(n19), .IN2(n28), .IN3(n23), .IN4(n29), .IN5(n30), .Q(B[7]) );
  AO222X1 U26 ( .IN1(n31), .IN2(n32), .IN3(n33), .IN4(n10), .IN5(n34), .IN6(
        n35), .Q(n30) );
  AO221X1 U27 ( .IN1(n19), .IN2(n36), .IN3(n23), .IN4(n37), .IN5(n38), .Q(B[6]) );
  AO222X1 U28 ( .IN1(n34), .IN2(n39), .IN3(n31), .IN4(n40), .IN5(n7), .IN6(n41), .Q(n38) );
  AO221X1 U29 ( .IN1(n19), .IN2(n42), .IN3(n23), .IN4(n20), .IN5(n43), .Q(B[5]) );
  AO222X1 U30 ( .IN1(n31), .IN2(n44), .IN3(n33), .IN4(n45), .IN5(n34), .IN6(
        n24), .Q(n43) );
  AO221X1 U31 ( .IN1(n19), .IN2(n46), .IN3(n23), .IN4(n25), .IN5(n47), .Q(B[4]) );
  AO222X1 U32 ( .IN1(n31), .IN2(n48), .IN3(n33), .IN4(n49), .IN5(n34), .IN6(
        n27), .Q(n47) );
  AND2X1 U33 ( .IN1(n41), .IN2(n8), .Q(n33) );
  NOR2X0 U34 ( .IN1(n50), .IN2(SH[7]), .QN(n41) );
  AND2X1 U35 ( .IN1(n21), .IN2(SH[2]), .Q(n31) );
  NOR2X0 U36 ( .IN1(SH[7]), .IN2(n51), .QN(B[3]) );
  OA222X1 U37 ( .IN1(n52), .IN2(n2), .IN3(n5), .IN4(n50), .IN5(n53), .IN6(n54), 
        .Q(n51) );
  OA221X1 U38 ( .IN1(n55), .IN2(n17), .IN3(n56), .IN4(n18), .IN5(n57), .Q(n53)
         );
  AOI22X1 U39 ( .IN1(n12), .IN2(A[5]), .IN3(n13), .IN4(A[6]), .QN(n57) );
  AOI222X1 U40 ( .IN1(n28), .IN2(n3), .IN3(n29), .IN4(n58), .IN5(n35), .IN6(
        n59), .QN(n52) );
  AO221X1 U41 ( .IN1(A[9]), .IN2(n12), .IN3(A[10]), .IN4(n13), .IN5(n60), .Q(
        n28) );
  AO22X1 U42 ( .IN1(A[7]), .IN2(n10), .IN3(A[8]), .IN4(n9), .Q(n60) );
  NOR2X0 U43 ( .IN1(SH[7]), .IN2(n61), .QN(B[2]) );
  OA222X1 U44 ( .IN1(n62), .IN2(n2), .IN3(n6), .IN4(n50), .IN5(n63), .IN6(n54), 
        .Q(n61) );
  OA221X1 U45 ( .IN1(n55), .IN2(n16), .IN3(n56), .IN4(n17), .IN5(n64), .Q(n63)
         );
  AOI22X1 U46 ( .IN1(n12), .IN2(A[4]), .IN3(n13), .IN4(A[5]), .QN(n64) );
  NAND2X0 U47 ( .IN1(n65), .IN2(n2), .QN(n50) );
  AOI222X1 U48 ( .IN1(n36), .IN2(n3), .IN3(n37), .IN4(n58), .IN5(n39), .IN6(
        n59), .QN(n62) );
  AO221X1 U49 ( .IN1(A[8]), .IN2(n12), .IN3(A[9]), .IN4(n13), .IN5(n67), .Q(
        n36) );
  AO22X1 U50 ( .IN1(A[6]), .IN2(n10), .IN3(A[7]), .IN4(n9), .Q(n67) );
  AND2X1 U51 ( .IN1(n10), .IN2(n19), .Q(B[23]) );
  NOR2X0 U52 ( .IN1(n68), .IN2(n69), .QN(B[22]) );
  AND2X1 U53 ( .IN1(n45), .IN2(n19), .Q(B[21]) );
  AND2X1 U54 ( .IN1(n49), .IN2(n19), .Q(B[20]) );
  OA21X1 U55 ( .IN1(n70), .IN2(n71), .IN3(n1), .Q(B[1]) );
  MUX21X1 U56 ( .IN1(n4), .IN2(n72), .S(n66), .Q(n71) );
  AO222X1 U57 ( .IN1(n59), .IN2(n24), .IN3(n58), .IN4(n20), .IN5(n3), .IN6(n42), .Q(n72) );
  AO221X1 U58 ( .IN1(A[7]), .IN2(n12), .IN3(A[8]), .IN4(n13), .IN5(n73), .Q(
        n42) );
  AO22X1 U59 ( .IN1(A[5]), .IN2(n10), .IN3(A[6]), .IN4(n9), .Q(n73) );
  AO221X1 U60 ( .IN1(A[11]), .IN2(n12), .IN3(A[12]), .IN4(n13), .IN5(n74), .Q(
        n20) );
  AO22X1 U61 ( .IN1(A[9]), .IN2(n10), .IN3(A[10]), .IN4(n9), .Q(n74) );
  NOR2X0 U62 ( .IN1(n76), .IN2(n54), .QN(n70) );
  OA221X1 U63 ( .IN1(n55), .IN2(n15), .IN3(n56), .IN4(n16), .IN5(n77), .Q(n76)
         );
  OA22X1 U64 ( .IN1(n78), .IN2(n17), .IN3(n79), .IN4(n18), .Q(n77) );
  NOR2X0 U65 ( .IN1(n5), .IN2(n69), .QN(B[19]) );
  NOR2X0 U66 ( .IN1(n6), .IN2(n69), .QN(B[18]) );
  NOR2X0 U67 ( .IN1(n81), .IN2(n75), .QN(B[17]) );
  NAND2X0 U68 ( .IN1(n65), .IN2(n22), .QN(n75) );
  MUX21X1 U69 ( .IN1(n45), .IN2(n44), .S(n8), .Q(n22) );
  NOR2X0 U70 ( .IN1(n81), .IN2(n83), .QN(B[16]) );
  AO222X1 U71 ( .IN1(n19), .IN2(n35), .IN3(n34), .IN4(n10), .IN5(n23), .IN6(
        n32), .Q(B[15]) );
  AO222X1 U72 ( .IN1(n7), .IN2(n21), .IN3(n19), .IN4(n39), .IN5(n23), .IN6(n40), .Q(B[14]) );
  NAND2X0 U73 ( .IN1(n84), .IN2(n8), .QN(n68) );
  AO222X1 U74 ( .IN1(n19), .IN2(n24), .IN3(n34), .IN4(n45), .IN5(n23), .IN6(
        n44), .Q(B[13]) );
  AO221X1 U75 ( .IN1(A[19]), .IN2(n12), .IN3(A[20]), .IN4(n13), .IN5(n85), .Q(
        n44) );
  AO22X1 U76 ( .IN1(A[17]), .IN2(n10), .IN3(A[18]), .IN4(n9), .Q(n85) );
  AO221X1 U77 ( .IN1(A[22]), .IN2(n9), .IN3(A[21]), .IN4(n14), .IN5(n12), .Q(
        n45) );
  AO221X1 U78 ( .IN1(A[15]), .IN2(n12), .IN3(A[16]), .IN4(n13), .IN5(n86), .Q(
        n24) );
  AO22X1 U79 ( .IN1(A[13]), .IN2(n10), .IN3(A[14]), .IN4(n9), .Q(n86) );
  AO222X1 U80 ( .IN1(n19), .IN2(n27), .IN3(n34), .IN4(n49), .IN5(n23), .IN6(
        n48), .Q(B[12]) );
  AND2X1 U81 ( .IN1(n21), .IN2(n8), .Q(n34) );
  AO222X1 U82 ( .IN1(n21), .IN2(n80), .IN3(n19), .IN4(n29), .IN5(n23), .IN6(
        n35), .Q(B[11]) );
  AO221X1 U83 ( .IN1(A[17]), .IN2(n12), .IN3(A[18]), .IN4(n13), .IN5(n87), .Q(
        n35) );
  AO22X1 U84 ( .IN1(A[15]), .IN2(n10), .IN3(A[16]), .IN4(n9), .Q(n87) );
  AO221X1 U85 ( .IN1(A[13]), .IN2(n12), .IN3(A[14]), .IN4(n13), .IN5(n88), .Q(
        n29) );
  AO22X1 U86 ( .IN1(A[11]), .IN2(n10), .IN3(A[12]), .IN4(n9), .Q(n88) );
  MUX21X1 U87 ( .IN1(n32), .IN2(n10), .S(SH[2]), .Q(n80) );
  AO221X1 U88 ( .IN1(n12), .IN2(A[21]), .IN3(n13), .IN4(A[22]), .IN5(n89), .Q(
        n32) );
  AO22X1 U89 ( .IN1(n10), .IN2(A[19]), .IN3(A[20]), .IN4(n9), .Q(n89) );
  AO222X1 U90 ( .IN1(n21), .IN2(n82), .IN3(n19), .IN4(n37), .IN5(n23), .IN6(
        n39), .Q(B[10]) );
  AO221X1 U91 ( .IN1(A[16]), .IN2(n12), .IN3(A[17]), .IN4(n13), .IN5(n90), .Q(
        n39) );
  AO22X1 U92 ( .IN1(A[14]), .IN2(n10), .IN3(A[15]), .IN4(n9), .Q(n90) );
  NOR2X0 U93 ( .IN1(n91), .IN2(n81), .QN(n23) );
  AO221X1 U94 ( .IN1(A[12]), .IN2(n12), .IN3(A[13]), .IN4(n13), .IN5(n92), .Q(
        n37) );
  AO22X1 U95 ( .IN1(A[10]), .IN2(n10), .IN3(A[11]), .IN4(n9), .Q(n92) );
  NOR2X0 U96 ( .IN1(n54), .IN2(SH[7]), .QN(n19) );
  MUX21X1 U97 ( .IN1(n40), .IN2(n84), .S(SH[2]), .Q(n82) );
  AO21X1 U98 ( .IN1(A[22]), .IN2(n11), .IN3(n9), .Q(n84) );
  AO221X1 U99 ( .IN1(A[20]), .IN2(n12), .IN3(n13), .IN4(A[21]), .IN5(n93), .Q(
        n40) );
  AO22X1 U100 ( .IN1(n10), .IN2(A[18]), .IN3(A[19]), .IN4(n9), .Q(n93) );
  NOR2X0 U101 ( .IN1(n81), .IN2(n65), .QN(n21) );
  NAND2X0 U102 ( .IN1(n66), .IN2(n1), .QN(n81) );
  NOR2X0 U103 ( .IN1(SH[7]), .IN2(n94), .QN(B[0]) );
  OA21X1 U104 ( .IN1(n95), .IN2(n54), .IN3(n96), .Q(n94) );
  MUX21X1 U105 ( .IN1(n83), .IN2(n97), .S(n66), .Q(n96) );
  AOI222X1 U106 ( .IN1(n46), .IN2(n3), .IN3(n25), .IN4(n58), .IN5(n27), .IN6(
        n59), .QN(n97) );
  NOR2X0 U107 ( .IN1(n8), .IN2(n65), .QN(n59) );
  AO221X1 U108 ( .IN1(A[14]), .IN2(n12), .IN3(A[15]), .IN4(n13), .IN5(n98), 
        .Q(n27) );
  AO22X1 U109 ( .IN1(A[12]), .IN2(n10), .IN3(A[13]), .IN4(n9), .Q(n98) );
  NOR2X0 U110 ( .IN1(n65), .IN2(SH[2]), .QN(n58) );
  AO221X1 U111 ( .IN1(A[10]), .IN2(n12), .IN3(A[11]), .IN4(n13), .IN5(n99), 
        .Q(n25) );
  AO22X1 U112 ( .IN1(A[8]), .IN2(n10), .IN3(A[9]), .IN4(n9), .Q(n99) );
  NAND2X0 U113 ( .IN1(n65), .IN2(SH[2]), .QN(n91) );
  AO221X1 U114 ( .IN1(A[6]), .IN2(n12), .IN3(A[7]), .IN4(n13), .IN5(n100), .Q(
        n46) );
  AO22X1 U115 ( .IN1(A[4]), .IN2(n10), .IN3(A[5]), .IN4(n9), .Q(n100) );
  NAND2X0 U116 ( .IN1(n65), .IN2(n26), .QN(n83) );
  MUX21X1 U117 ( .IN1(n49), .IN2(n48), .S(n8), .Q(n26) );
  AO221X1 U118 ( .IN1(A[18]), .IN2(n12), .IN3(n13), .IN4(A[19]), .IN5(n101), 
        .Q(n48) );
  AO22X1 U119 ( .IN1(A[16]), .IN2(n10), .IN3(A[17]), .IN4(n9), .Q(n101) );
  AO221X1 U120 ( .IN1(A[21]), .IN2(SH[0]), .IN3(A[22]), .IN4(SH[1]), .IN5(n102), .Q(n49) );
  AO21X1 U121 ( .IN1(n10), .IN2(A[20]), .IN3(n13), .Q(n102) );
  NAND3X0 U122 ( .IN1(n66), .IN2(n8), .IN3(n65), .QN(n54) );
  NOR2X0 U123 ( .IN1(SH[4]), .IN2(n103), .QN(n66) );
  OR2X1 U124 ( .IN1(SH[5]), .IN2(SH[6]), .Q(n103) );
  OA221X1 U125 ( .IN1(n79), .IN2(n17), .IN3(n78), .IN4(n16), .IN5(n104), .Q(
        n95) );
  AOI22X1 U126 ( .IN1(A[1]), .IN2(n9), .IN3(A[0]), .IN4(n10), .QN(n104) );
  NAND2X0 U127 ( .IN1(n14), .IN2(n11), .QN(n55) );
  NAND2X0 U128 ( .IN1(SH[0]), .IN2(n11), .QN(n56) );
  NAND2X0 U129 ( .IN1(SH[1]), .IN2(n14), .QN(n78) );
  NAND2X0 U130 ( .IN1(SH[0]), .IN2(SH[1]), .QN(n79) );
endmodule


module fpalu_add1_DW01_sub_25 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8;
  wire   [8:0] carry;

  FADDX1 U2_6 ( .A(A[6]), .B(n7), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FADDX1 U2_5 ( .A(A[5]), .B(n6), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FADDX1 U2_4 ( .A(A[4]), .B(n5), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FADDX1 U2_3 ( .A(A[3]), .B(n4), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  FADDX1 U2_2 ( .A(A[2]), .B(n3), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  FADDX1 U2_1 ( .A(A[1]), .B(n2), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  XOR3X1 U2_7 ( .IN1(A[7]), .IN2(n8), .IN3(carry[7]), .Q(DIFF[7]) );
  NAND2X1 U1 ( .IN1(n1), .IN2(B[0]), .QN(carry[1]) );
  INVX0 U2 ( .INP(B[1]), .ZN(n2) );
  INVX0 U3 ( .INP(A[0]), .ZN(n1) );
  INVX0 U4 ( .INP(B[2]), .ZN(n3) );
  INVX0 U5 ( .INP(B[5]), .ZN(n6) );
  INVX0 U6 ( .INP(B[6]), .ZN(n7) );
  INVX0 U7 ( .INP(B[4]), .ZN(n5) );
  INVX0 U8 ( .INP(B[3]), .ZN(n4) );
  INVX0 U9 ( .INP(B[7]), .ZN(n8) );
  XOR2X1 U10 ( .IN1(B[0]), .IN2(A[0]), .Q(DIFF[0]) );
endmodule


module fpalu_add1 ( a_in, b_in, sum, overflow );
  input [31:0] a_in;
  input [31:0] b_in;
  output [31:0] sum;
  output overflow;
  wire   sum_31, N54, N59, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72,
         N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86,
         N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N117,
         N118, N119, N120, N121, N122, N123, N124, N125, N126, N127, N128,
         N129, N130, N131, N132, N133, N134, N135, N136, N137, N138, N139,
         N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161,
         N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172,
         N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183,
         N184, N185, N186, N187, N188, N213, N214, N215, N216, N217, N218,
         N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229,
         N230, N231, N232, N233, N234, N235, N236, N237, N241, N242, N243,
         N244, N245, N246, N247, N248, N249, N250, N251, N252, N253, N254,
         N255, N256, N257, N258, N259, N260, N261, N262, N263, N264, N290,
         N291, N292, N293, N294, N295, N296, N297, N368, N369, N370, N371,
         N372, N373, N374, N375, N436, N438, N439, N440, N441, N442, N443,
         N549, N550, N551, N552, N553, N554, N555, N662, N664, N665, N666,
         N667, N668, N775, N776, N777, N778, N779, N780, N781, N889, N890,
         N891, N892, N893, N894, N1001, N1002, N1003, N1004, N1005, N1006,
         N1007, N1116, N1118, N1119, N1120, N1121, N1230, N1231, N1232, N1233,
         N1234, N1235, N1236, N1346, N1347, N1348, N1349, N1350, N1351, N1460,
         N1461, N1462, N1463, N1464, N1465, N1466, N1577, N1578, N1579, N1580,
         N1581, N1690, N1691, N1692, N1693, N1694, N1695, N1696, N1806, N1807,
         N1808, N1809, N1810, N1811, N1920, N1921, N1922, N1923, N1924, N1925,
         N1926, N2037, N2039, N2040, N2041, N2150, N2151, N2152, N2153, N2154,
         N2155, N2156, N2266, N2267, N2268, N2269, N2270, N2271, N2380, N2381,
         N2382, N2383, N2384, N2385, N2386, N2497, N2498, N2499, N2500, N2501,
         N2610, N2611, N2612, N2613, N2614, N2615, N2616, N2726, N2727, N2728,
         N2729, N2730, N2731, N2764, N2765, N2766, N2767, N2768, N2802, N2803,
         N2804, N2805, N2806, N2807, N2808, N2809, N2810, N2811,
         \sub_114_I23/carry[7] , \sub_114_I23/carry[6] ,
         \sub_114_I23/carry[5] , \sub_114_I23/carry[4] ,
         \sub_114_I23/carry[3] , \sub_114_I22/carry[2] ,
         \sub_114_I22/carry[3] , \sub_114_I22/carry[4] ,
         \sub_114_I22/carry[5] , \sub_114_I22/carry[6] ,
         \sub_114_I22/carry[7] , \sub_114_I21/carry[7] ,
         \sub_114_I21/carry[6] , \sub_114_I21/carry[5] ,
         \sub_114_I21/carry[4] , \sub_114_I20/carry[2] ,
         \sub_114_I20/carry[3] , \sub_114_I20/carry[4] ,
         \sub_114_I20/carry[5] , \sub_114_I20/carry[6] ,
         \sub_114_I20/carry[7] , \sub_114_I19/carry[7] ,
         \sub_114_I19/carry[6] , \sub_114_I19/carry[5] ,
         \sub_114_I19/carry[4] , \sub_114_I19/carry[3] ,
         \sub_114_I18/carry[2] , \sub_114_I18/carry[3] ,
         \sub_114_I18/carry[4] , \sub_114_I18/carry[5] ,
         \sub_114_I18/carry[6] , \sub_114_I18/carry[7] ,
         \sub_114_I17/carry[7] , \sub_114_I17/carry[6] ,
         \sub_114_I16/carry[2] , \sub_114_I16/carry[3] ,
         \sub_114_I16/carry[4] , \sub_114_I16/carry[5] ,
         \sub_114_I16/carry[6] , \sub_114_I16/carry[7] ,
         \sub_114_I15/carry[7] , \sub_114_I15/carry[6] ,
         \sub_114_I15/carry[5] , \sub_114_I15/carry[4] ,
         \sub_114_I15/carry[3] , \sub_114_I14/carry[2] ,
         \sub_114_I14/carry[3] , \sub_114_I14/carry[4] ,
         \sub_114_I14/carry[5] , \sub_114_I14/carry[6] ,
         \sub_114_I14/carry[7] , \sub_114_I13/carry[7] ,
         \sub_114_I13/carry[6] , \sub_114_I13/carry[5] ,
         \sub_114_I13/carry[4] , \sub_114_I12/carry[2] ,
         \sub_114_I12/carry[3] , \sub_114_I12/carry[4] ,
         \sub_114_I12/carry[5] , \sub_114_I12/carry[6] ,
         \sub_114_I12/carry[7] , \sub_114_I11/carry[7] ,
         \sub_114_I11/carry[6] , \sub_114_I11/carry[5] ,
         \sub_114_I11/carry[4] , \sub_114_I11/carry[3] ,
         \sub_114_I10/carry[2] , \sub_114_I10/carry[3] ,
         \sub_114_I10/carry[4] , \sub_114_I10/carry[5] ,
         \sub_114_I10/carry[6] , \sub_114_I10/carry[7] , \sub_114_I9/carry[7] ,
         \sub_114_I9/carry[6] , \sub_114_I9/carry[5] , \sub_114_I8/carry[2] ,
         \sub_114_I8/carry[3] , \sub_114_I8/carry[4] , \sub_114_I8/carry[5] ,
         \sub_114_I8/carry[6] , \sub_114_I8/carry[7] , \sub_114_I7/carry[7] ,
         \sub_114_I7/carry[6] , \sub_114_I7/carry[5] , \sub_114_I7/carry[4] ,
         \sub_114_I7/carry[3] , \sub_114_I6/carry[2] , \sub_114_I6/carry[3] ,
         \sub_114_I6/carry[4] , \sub_114_I6/carry[5] , \sub_114_I6/carry[6] ,
         \sub_114_I6/carry[7] , \sub_114_I5/carry[7] , \sub_114_I5/carry[6] ,
         \sub_114_I5/carry[5] , \sub_114_I5/carry[4] , \sub_114_I4/carry[2] ,
         \sub_114_I4/carry[3] , \sub_114_I4/carry[4] , \sub_114_I4/carry[5] ,
         \sub_114_I4/carry[6] , \sub_114_I4/carry[7] , \sub_114_I3/carry[7] ,
         \sub_114_I3/carry[6] , \sub_114_I3/carry[5] , \sub_114_I3/carry[4] ,
         \sub_114_I3/carry[3] , \sub_114_I2_aco/carry[7] ,
         \sub_114_I2_aco/carry[6] , \sub_114_I2_aco/carry[5] ,
         \sub_114_I2_aco/carry[4] , \sub_114_I2_aco/carry[3] ,
         \sub_114_I2_aco/carry[2] , \sub_114_I2_aco/carry[1] ,
         \sub_114_I2_aco/B[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610;
  wire   [31:0] a;
  wire   [31:0] b;
  wire   [23:0] bsig;
  wire   [7:0] shift;
  wire   [23:0] asig1;
  wire   [23:0] bsig1;
  wire   [7:0] sumexp;
  wire   [31:0] x;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign sum[31] = sum_31;
  assign sum[30] = sumexp[7];
  assign sum[29] = sumexp[6];
  assign sum[28] = sumexp[5];
  assign sum[27] = sumexp[4];
  assign sum[26] = sumexp[3];
  assign sum[25] = sumexp[2];
  assign sum[24] = sumexp[1];
  assign sum[23] = sumexp[0];

  LATCHX1 \asig1_reg[23]  ( .CLK(a[31]), .D(N86), .Q(asig1[23]) );
  LATCHX1 \asig1_reg[22]  ( .CLK(a[31]), .D(N85), .Q(asig1[22]) );
  LATCHX1 \asig1_reg[21]  ( .CLK(a[31]), .D(N84), .Q(asig1[21]) );
  LATCHX1 \asig1_reg[20]  ( .CLK(a[31]), .D(N83), .Q(asig1[20]) );
  LATCHX1 \asig1_reg[19]  ( .CLK(a[31]), .D(N82), .Q(asig1[19]) );
  LATCHX1 \asig1_reg[18]  ( .CLK(n30), .D(N81), .Q(asig1[18]) );
  LATCHX1 \asig1_reg[17]  ( .CLK(n30), .D(N80), .Q(asig1[17]) );
  LATCHX1 \asig1_reg[16]  ( .CLK(n30), .D(N79), .Q(asig1[16]) );
  LATCHX1 \asig1_reg[15]  ( .CLK(n30), .D(N78), .Q(asig1[15]) );
  LATCHX1 \asig1_reg[14]  ( .CLK(n30), .D(N77), .Q(asig1[14]) );
  LATCHX1 \asig1_reg[13]  ( .CLK(n30), .D(N76), .Q(asig1[13]) );
  LATCHX1 \asig1_reg[12]  ( .CLK(n30), .D(N75), .Q(asig1[12]) );
  LATCHX1 \asig1_reg[11]  ( .CLK(n30), .D(N74), .Q(asig1[11]) );
  LATCHX1 \asig1_reg[10]  ( .CLK(n30), .D(N73), .Q(asig1[10]) );
  LATCHX1 \asig1_reg[9]  ( .CLK(n30), .D(N72), .Q(asig1[9]) );
  LATCHX1 \asig1_reg[8]  ( .CLK(n30), .D(N71), .Q(asig1[8]) );
  LATCHX1 \asig1_reg[7]  ( .CLK(n30), .D(N70), .Q(asig1[7]) );
  LATCHX1 \asig1_reg[6]  ( .CLK(n30), .D(N69), .Q(asig1[6]) );
  LATCHX1 \asig1_reg[5]  ( .CLK(n30), .D(N68), .Q(asig1[5]) );
  LATCHX1 \asig1_reg[4]  ( .CLK(n30), .D(N67), .Q(asig1[4]) );
  LATCHX1 \asig1_reg[3]  ( .CLK(n30), .D(N66), .Q(asig1[3]) );
  LATCHX1 \asig1_reg[2]  ( .CLK(n30), .D(N65), .Q(asig1[2]) );
  LATCHX1 \asig1_reg[1]  ( .CLK(n30), .D(N64), .Q(asig1[1]) );
  LATCHX1 \asig1_reg[0]  ( .CLK(n30), .D(N63), .Q(asig1[0]) );
  LATCHX1 \bsig1_reg[23]  ( .CLK(b[31]), .D(N110), .Q(bsig1[23]) );
  LATCHX1 \bsig1_reg[22]  ( .CLK(b[31]), .D(N109), .Q(bsig1[22]) );
  LATCHX1 \bsig1_reg[21]  ( .CLK(b[31]), .D(N108), .Q(bsig1[21]) );
  LATCHX1 \bsig1_reg[20]  ( .CLK(b[31]), .D(N107), .Q(bsig1[20]) );
  LATCHX1 \bsig1_reg[19]  ( .CLK(b[31]), .D(N106), .Q(bsig1[19]) );
  LATCHX1 \bsig1_reg[18]  ( .CLK(n24), .D(N105), .Q(bsig1[18]) );
  LATCHX1 \bsig1_reg[17]  ( .CLK(n24), .D(N104), .Q(bsig1[17]) );
  LATCHX1 \bsig1_reg[16]  ( .CLK(n24), .D(N103), .Q(bsig1[16]) );
  LATCHX1 \bsig1_reg[15]  ( .CLK(n24), .D(N102), .Q(bsig1[15]) );
  LATCHX1 \bsig1_reg[14]  ( .CLK(n24), .D(N101), .Q(bsig1[14]) );
  LATCHX1 \bsig1_reg[13]  ( .CLK(n24), .D(N100), .Q(bsig1[13]) );
  LATCHX1 \bsig1_reg[12]  ( .CLK(n24), .D(N99), .Q(bsig1[12]) );
  LATCHX1 \bsig1_reg[11]  ( .CLK(n24), .D(N98), .Q(bsig1[11]) );
  LATCHX1 \bsig1_reg[10]  ( .CLK(n24), .D(N97), .Q(bsig1[10]) );
  LATCHX1 \bsig1_reg[9]  ( .CLK(n24), .D(N96), .Q(bsig1[9]) );
  LATCHX1 \bsig1_reg[8]  ( .CLK(n24), .D(N95), .Q(bsig1[8]) );
  LATCHX1 \bsig1_reg[7]  ( .CLK(n24), .D(N94), .Q(bsig1[7]) );
  LATCHX1 \bsig1_reg[6]  ( .CLK(n24), .D(N93), .Q(bsig1[6]) );
  LATCHX1 \bsig1_reg[5]  ( .CLK(n24), .D(N92), .Q(bsig1[5]) );
  LATCHX1 \bsig1_reg[4]  ( .CLK(n24), .D(N91), .Q(bsig1[4]) );
  LATCHX1 \bsig1_reg[3]  ( .CLK(n24), .D(N90), .Q(bsig1[3]) );
  LATCHX1 \bsig1_reg[2]  ( .CLK(n24), .D(N89), .Q(bsig1[2]) );
  LATCHX1 \bsig1_reg[1]  ( .CLK(n24), .D(N88), .Q(bsig1[1]) );
  LATCHX1 \bsig1_reg[0]  ( .CLK(n24), .D(N87), .Q(bsig1[0]) );
  LATCHX1 \x_reg[3]  ( .CLK(N2811), .D(N2767), .Q(x[3]) );
  LATCHX1 \x_reg[0]  ( .CLK(N2811), .D(N2764), .Q(x[0]) );
  LATCHX1 \x_reg[4]  ( .CLK(N2811), .D(N2768), .Q(x[4]) );
  LATCHX1 \x_reg[2]  ( .CLK(N2811), .D(N2766), .Q(x[2]) );
  LATCHX1 \x_reg[1]  ( .CLK(N2811), .D(N2765), .Q(x[1]) );
  LATCHX1 \sumexp_reg[7]  ( .CLK(N2802), .D(N2810), .Q(sumexp[7]) );
  LATCHX1 \sumexp_reg[6]  ( .CLK(N2802), .D(N2809), .Q(sumexp[6]) );
  LATCHX1 \sumexp_reg[5]  ( .CLK(N2802), .D(N2808), .Q(sumexp[5]) );
  LATCHX1 \sumexp_reg[4]  ( .CLK(N2802), .D(N2807), .Q(sumexp[4]) );
  LATCHX1 \sumexp_reg[3]  ( .CLK(N2802), .D(N2806), .Q(sumexp[3]) );
  LATCHX1 \sumexp_reg[2]  ( .CLK(N2802), .D(N2805), .Q(sumexp[2]) );
  LATCHX1 \sumexp_reg[1]  ( .CLK(N2802), .D(N2804), .Q(sumexp[1]) );
  LATCHX1 \sumexp_reg[0]  ( .CLK(N2802), .D(N2803), .Q(sumexp[0]) );
  fpalu_add1_DW01_inc_0 add_83 ( .A({a[30:29], n8, n7, n3, n20, n5, N436}), 
        .SUM({N297, N296, N295, N294, N293, N292, N291, N290}) );
  fpalu_add1_DW01_sub_22 sub_77 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({N236, N235, N234, N233, N232, N231, 
        N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, 
        N218, N217, N216, N215, N214, N213}), .CI(1'b0), .DIFF({N264, N263, 
        N262, N261, N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, 
        N250, N249, N248, N247, N246, N245, N244, N243, N242, N241}) );
  fpalu_add1_DW01_add_0 add_69 ( .A(asig1), .B(bsig), .CI(1'b0), .SUM({N188, 
        N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, 
        N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, N165}) );
  fpalu_add1_DW01_add_1 add_68 ( .A({1'b1, a[22:0]}), .B(bsig1), .CI(1'b0), 
        .SUM({N164, N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, 
        N153, N152, N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, 
        N141}) );
  fpalu_add1_DW01_sub_23 sub_61_S2 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({1'b0, bsig}), .CI(1'b0), .DIFF({SYNOPSYS_UNCONNECTED__0, N110, N109, N108, N107, N106, N105, N104, 
        N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, 
        N90, N89, N88, N87}) );
  fpalu_add1_DW01_sub_24 sub_60_S2 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({1'b0, 1'b1, a[22:0]}), 
        .CI(1'b0), .DIFF({SYNOPSYS_UNCONNECTED__1, N86, N85, N84, N83, N82, 
        N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, 
        N67, N66, N65, N64, N63}) );
  fpalu_add1_DW01_add_2 r357 ( .A({1'b1, a[22:0]}), .B(bsig), .CI(1'b0), .SUM(
        {N140, N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, 
        N129, N128, N127, N126, N125, N124, N123, N122, N121, N120, N119, N118, 
        N117}) );
  fpalu_add1_DW01_cmp6_0 r354 ( .A({1'b0, 1'b0, 1'b1, a[22:0]}), .B({1'b0, 
        1'b0, bsig}), .TC(1'b0), .LT(N237), .GT(N59) );
  fpalu_add1_DW_rash_0 srl_47 ( .A({1'b1, b[22:0]}), .DATA_TC(1'b0), .SH(shift), .SH_TC(1'b0), .B(bsig) );
  fpalu_add1_DW01_sub_25 sub_46 ( .A({a[30:29], n8, n6, n2, n20, n4, N436}), 
        .B(b[30:23]), .CI(1'b0), .DIFF(shift) );
  AND4X1 U3 ( .IN1(n68), .IN2(n81), .IN3(n82), .IN4(n83), .Q(n1) );
  NOR2X0 U4 ( .IN1(n25), .IN2(a[31]), .QN(n608) );
  AO21X1 U5 ( .IN1(n86), .IN2(n65), .IN3(n1), .Q(sum[6]) );
  NOR2X0 U6 ( .IN1(n31), .IN2(b[31]), .QN(n607) );
  XOR2X1 U7 ( .IN1(\sub_114_I18/carry[2] ), .IN2(n21), .Q(N2151) );
  AO221X1 U8 ( .IN1(N372), .IN2(n348), .IN3(N440), .IN4(n177), .IN5(n391), .Q(
        n388) );
  XNOR2X1 U9 ( .IN1(n21), .IN2(\sub_114_I22/carry[2] ), .Q(N2611) );
  XNOR2X1 U10 ( .IN1(\sub_114_I18/carry[6] ), .IN2(a[29]), .Q(N2155) );
  AO22X1 U11 ( .IN1(n176), .IN2(n65), .IN3(n241), .IN4(n76), .Q(sum[17]) );
  AND3X1 U12 ( .IN1(n507), .IN2(n531), .IN3(n155), .Q(n516) );
  XOR2X1 U13 ( .IN1(\sub_114_I20/carry[2] ), .IN2(n21), .Q(N2381) );
  OR2X1 U14 ( .IN1(a[29]), .IN2(\sub_114_I20/carry[6] ), .Q(
        \sub_114_I20/carry[7] ) );
  OA21X1 U15 ( .IN1(n324), .IN2(n322), .IN3(n13), .Q(N2811) );
  INVX0 U16 ( .INP(n65), .ZN(n13) );
  INVX0 U17 ( .INP(n121), .ZN(\sub_114_I2_aco/B[0] ) );
  NBUFFX2 U18 ( .INP(n457), .Z(n15) );
  NBUFFX2 U19 ( .INP(n177), .Z(n14) );
  NBUFFX2 U20 ( .INP(n607), .Z(n16) );
  NBUFFX4 U21 ( .INP(a[28]), .Z(n9) );
  AND2X1 U22 ( .IN1(n145), .IN2(n121), .Q(n175) );
  NBUFFX4 U23 ( .INP(a[29]), .Z(n11) );
  NBUFFX4 U24 ( .INP(a[29]), .Z(n10) );
  NBUFFX2 U25 ( .INP(n608), .Z(n17) );
  NBUFFX4 U26 ( .INP(a[27]), .Z(n7) );
  NBUFFX4 U27 ( .INP(N2037), .Z(n3) );
  NBUFFX4 U28 ( .INP(N662), .Z(n5) );
  NBUFFX2 U29 ( .INP(a[28]), .Z(n8) );
  NBUFFX2 U30 ( .INP(n610), .Z(n18) );
  NBUFFX2 U31 ( .INP(a[27]), .Z(n6) );
  NBUFFX2 U32 ( .INP(N662), .Z(n4) );
  NBUFFX2 U33 ( .INP(N2037), .Z(n2) );
  NAND3X0 U34 ( .IN1(n529), .IN2(n459), .IN3(n508), .QN(n152) );
  NAND3X0 U35 ( .IN1(n582), .IN2(n540), .IN3(n550), .QN(n185) );
  AND2X1 U36 ( .IN1(n443), .IN2(n83), .Q(n339) );
  NAND3X0 U37 ( .IN1(n539), .IN2(n540), .IN3(n541), .QN(n151) );
  NBUFFX2 U38 ( .INP(N54), .Z(n36) );
  NBUFFX2 U39 ( .INP(N54), .Z(n32) );
  NBUFFX2 U40 ( .INP(N54), .Z(n33) );
  NBUFFX2 U41 ( .INP(N54), .Z(n34) );
  NBUFFX2 U42 ( .INP(N54), .Z(n35) );
  NAND3X0 U43 ( .IN1(n583), .IN2(n540), .IN3(n477), .QN(n182) );
  NAND3X0 U44 ( .IN1(n554), .IN2(n540), .IN3(n555), .QN(n205) );
  NAND3X0 U45 ( .IN1(n528), .IN2(n459), .IN3(n518), .QN(n83) );
  NOR4X0 U46 ( .IN1(x[1]), .IN2(x[0]), .IN3(x[2]), .IN4(n609), .QN(n510) );
  INVX0 U47 ( .INP(a_in[30]), .ZN(n62) );
  INVX0 U48 ( .INP(a[27]), .ZN(n26) );
  INVX0 U49 ( .INP(N1116), .ZN(n21) );
  INVX0 U50 ( .INP(b_in[23]), .ZN(n55) );
  INVX0 U51 ( .INP(a[28]), .ZN(n27) );
  INVX0 U52 ( .INP(N662), .ZN(n22) );
  INVX0 U53 ( .INP(N436), .ZN(n23) );
  INVX0 U54 ( .INP(N2037), .ZN(n19) );
  INVX0 U55 ( .INP(b[31]), .ZN(n25) );
  INVX0 U56 ( .INP(a_in[25]), .ZN(n57) );
  INVX0 U57 ( .INP(a[30]), .ZN(n29) );
  INVX0 U58 ( .INP(a[29]), .ZN(n28) );
  INVX0 U59 ( .INP(a_in[28]), .ZN(n60) );
  INVX0 U60 ( .INP(a_in[26]), .ZN(n58) );
  INVX0 U61 ( .INP(a_in[27]), .ZN(n59) );
  INVX0 U62 ( .INP(a_in[24]), .ZN(n56) );
  INVX0 U63 ( .INP(a_in[29]), .ZN(n61) );
  INVX0 U64 ( .INP(n13), .ZN(n12) );
  INVX0 U65 ( .INP(n21), .ZN(n20) );
  INVX0 U66 ( .INP(n25), .ZN(n24) );
  INVX0 U67 ( .INP(n31), .ZN(n30) );
  INVX0 U68 ( .INP(a[31]), .ZN(n31) );
  XNOR2X1 U69 ( .IN1(a[30]), .IN2(\sub_114_I23/carry[7] ), .Q(N2731) );
  OR2X1 U70 ( .IN1(a[29]), .IN2(\sub_114_I23/carry[6] ), .Q(
        \sub_114_I23/carry[7] ) );
  XNOR2X1 U71 ( .IN1(\sub_114_I23/carry[6] ), .IN2(n11), .Q(N2730) );
  OR2X1 U72 ( .IN1(a[28]), .IN2(\sub_114_I23/carry[5] ), .Q(
        \sub_114_I23/carry[6] ) );
  XNOR2X1 U73 ( .IN1(\sub_114_I23/carry[5] ), .IN2(n9), .Q(N2729) );
  AND2X1 U74 ( .IN1(\sub_114_I23/carry[4] ), .IN2(n6), .Q(
        \sub_114_I23/carry[5] ) );
  XOR2X1 U84 ( .IN1(n7), .IN2(\sub_114_I23/carry[4] ), .Q(N2728) );
  OR2X1 U85 ( .IN1(n2), .IN2(\sub_114_I23/carry[3] ), .Q(
        \sub_114_I23/carry[4] ) );
  XNOR2X1 U86 ( .IN1(\sub_114_I23/carry[3] ), .IN2(N2037), .Q(N2727) );
  AND2X1 U87 ( .IN1(n4), .IN2(N1116), .Q(\sub_114_I23/carry[3] ) );
  XOR2X1 U88 ( .IN1(n20), .IN2(n5), .Q(N2726) );
  XNOR2X1 U89 ( .IN1(a[30]), .IN2(\sub_114_I22/carry[7] ), .Q(N2616) );
  OR2X1 U90 ( .IN1(a[29]), .IN2(\sub_114_I22/carry[6] ), .Q(
        \sub_114_I22/carry[7] ) );
  XNOR2X1 U91 ( .IN1(\sub_114_I22/carry[6] ), .IN2(n11), .Q(N2615) );
  OR2X1 U92 ( .IN1(a[28]), .IN2(\sub_114_I22/carry[5] ), .Q(
        \sub_114_I22/carry[6] ) );
  XNOR2X1 U93 ( .IN1(\sub_114_I22/carry[5] ), .IN2(n9), .Q(N2614) );
  AND2X1 U94 ( .IN1(\sub_114_I22/carry[4] ), .IN2(a[27]), .Q(
        \sub_114_I22/carry[5] ) );
  XOR2X1 U95 ( .IN1(n7), .IN2(\sub_114_I22/carry[4] ), .Q(N2613) );
  OR2X1 U96 ( .IN1(N2037), .IN2(\sub_114_I22/carry[3] ), .Q(
        \sub_114_I22/carry[4] ) );
  XNOR2X1 U97 ( .IN1(\sub_114_I22/carry[3] ), .IN2(n3), .Q(N2612) );
  AND2X1 U98 ( .IN1(\sub_114_I22/carry[2] ), .IN2(N1116), .Q(
        \sub_114_I22/carry[3] ) );
  OR2X1 U99 ( .IN1(N662), .IN2(N436), .Q(\sub_114_I22/carry[2] ) );
  XNOR2X1 U100 ( .IN1(N436), .IN2(n5), .Q(N2610) );
  XNOR2X1 U101 ( .IN1(a[30]), .IN2(\sub_114_I19/carry[7] ), .Q(N2271) );
  OR2X1 U102 ( .IN1(a[29]), .IN2(\sub_114_I19/carry[6] ), .Q(
        \sub_114_I19/carry[7] ) );
  XNOR2X1 U103 ( .IN1(\sub_114_I19/carry[6] ), .IN2(n11), .Q(N2270) );
  OR2X1 U104 ( .IN1(a[28]), .IN2(\sub_114_I19/carry[5] ), .Q(
        \sub_114_I19/carry[6] ) );
  XNOR2X1 U105 ( .IN1(\sub_114_I19/carry[5] ), .IN2(n9), .Q(N2269) );
  AND2X1 U106 ( .IN1(\sub_114_I19/carry[4] ), .IN2(n6), .Q(
        \sub_114_I19/carry[5] ) );
  XOR2X1 U107 ( .IN1(n7), .IN2(\sub_114_I19/carry[4] ), .Q(N2268) );
  OR2X1 U108 ( .IN1(N2037), .IN2(\sub_114_I19/carry[3] ), .Q(
        \sub_114_I19/carry[4] ) );
  XNOR2X1 U109 ( .IN1(\sub_114_I19/carry[3] ), .IN2(n3), .Q(N2267) );
  OR2X1 U110 ( .IN1(N1116), .IN2(n5), .Q(\sub_114_I19/carry[3] ) );
  XNOR2X1 U111 ( .IN1(n4), .IN2(n20), .Q(N2266) );
  XNOR2X1 U112 ( .IN1(a[30]), .IN2(\sub_114_I17/carry[7] ), .Q(N2041) );
  OR2X1 U113 ( .IN1(a[29]), .IN2(\sub_114_I17/carry[6] ), .Q(
        \sub_114_I17/carry[7] ) );
  XNOR2X1 U114 ( .IN1(\sub_114_I17/carry[6] ), .IN2(n11), .Q(N2040) );
  OR2X1 U115 ( .IN1(a[28]), .IN2(n6), .Q(\sub_114_I17/carry[6] ) );
  XNOR2X1 U116 ( .IN1(a[27]), .IN2(n9), .Q(N2039) );
  XNOR2X1 U117 ( .IN1(a[30]), .IN2(\sub_114_I21/carry[7] ), .Q(N2501) );
  OR2X1 U118 ( .IN1(a[29]), .IN2(\sub_114_I21/carry[6] ), .Q(
        \sub_114_I21/carry[7] ) );
  XNOR2X1 U119 ( .IN1(\sub_114_I21/carry[6] ), .IN2(n11), .Q(N2500) );
  OR2X1 U120 ( .IN1(a[28]), .IN2(\sub_114_I21/carry[5] ), .Q(
        \sub_114_I21/carry[6] ) );
  XNOR2X1 U121 ( .IN1(\sub_114_I21/carry[5] ), .IN2(n9), .Q(N2499) );
  AND2X1 U122 ( .IN1(\sub_114_I21/carry[4] ), .IN2(a[27]), .Q(
        \sub_114_I21/carry[5] ) );
  XOR2X1 U123 ( .IN1(n6), .IN2(\sub_114_I21/carry[4] ), .Q(N2498) );
  OR2X1 U124 ( .IN1(N2037), .IN2(N1116), .Q(\sub_114_I21/carry[4] ) );
  XNOR2X1 U125 ( .IN1(N1116), .IN2(N2037), .Q(N2497) );
  XNOR2X1 U126 ( .IN1(a[30]), .IN2(\sub_114_I18/carry[7] ), .Q(N2156) );
  OR2X1 U127 ( .IN1(n10), .IN2(\sub_114_I18/carry[6] ), .Q(
        \sub_114_I18/carry[7] ) );
  OR2X1 U128 ( .IN1(a[28]), .IN2(\sub_114_I18/carry[5] ), .Q(
        \sub_114_I18/carry[6] ) );
  XNOR2X1 U129 ( .IN1(\sub_114_I18/carry[5] ), .IN2(n9), .Q(N2154) );
  AND2X1 U130 ( .IN1(\sub_114_I18/carry[4] ), .IN2(n6), .Q(
        \sub_114_I18/carry[5] ) );
  XOR2X1 U131 ( .IN1(n7), .IN2(\sub_114_I18/carry[4] ), .Q(N2153) );
  OR2X1 U132 ( .IN1(n2), .IN2(\sub_114_I18/carry[3] ), .Q(
        \sub_114_I18/carry[4] ) );
  XNOR2X1 U133 ( .IN1(\sub_114_I18/carry[3] ), .IN2(N2037), .Q(N2152) );
  OR2X1 U134 ( .IN1(N1116), .IN2(\sub_114_I18/carry[2] ), .Q(
        \sub_114_I18/carry[3] ) );
  OR2X1 U135 ( .IN1(N662), .IN2(N436), .Q(\sub_114_I18/carry[2] ) );
  XNOR2X1 U136 ( .IN1(N436), .IN2(n5), .Q(N2150) );
  XNOR2X1 U137 ( .IN1(a[30]), .IN2(\sub_114_I20/carry[7] ), .Q(N2386) );
  XNOR2X1 U138 ( .IN1(\sub_114_I20/carry[6] ), .IN2(n11), .Q(N2385) );
  OR2X1 U139 ( .IN1(n9), .IN2(\sub_114_I20/carry[5] ), .Q(
        \sub_114_I20/carry[6] ) );
  XNOR2X1 U140 ( .IN1(\sub_114_I20/carry[5] ), .IN2(n9), .Q(N2384) );
  AND2X1 U141 ( .IN1(\sub_114_I20/carry[4] ), .IN2(a[27]), .Q(
        \sub_114_I20/carry[5] ) );
  XOR2X1 U142 ( .IN1(n6), .IN2(\sub_114_I20/carry[4] ), .Q(N2383) );
  OR2X1 U143 ( .IN1(n2), .IN2(\sub_114_I20/carry[3] ), .Q(
        \sub_114_I20/carry[4] ) );
  XNOR2X1 U144 ( .IN1(\sub_114_I20/carry[3] ), .IN2(n3), .Q(N2382) );
  OR2X1 U145 ( .IN1(N1116), .IN2(\sub_114_I20/carry[2] ), .Q(
        \sub_114_I20/carry[3] ) );
  AND2X1 U146 ( .IN1(N436), .IN2(n4), .Q(\sub_114_I20/carry[2] ) );
  XOR2X1 U147 ( .IN1(n5), .IN2(N436), .Q(N2380) );
  XNOR2X1 U148 ( .IN1(a[30]), .IN2(\sub_114_I13/carry[7] ), .Q(N1581) );
  OR2X1 U149 ( .IN1(n10), .IN2(\sub_114_I13/carry[6] ), .Q(
        \sub_114_I13/carry[7] ) );
  XNOR2X1 U150 ( .IN1(\sub_114_I13/carry[6] ), .IN2(n11), .Q(N1580) );
  OR2X1 U151 ( .IN1(n9), .IN2(\sub_114_I13/carry[5] ), .Q(
        \sub_114_I13/carry[6] ) );
  XNOR2X1 U152 ( .IN1(\sub_114_I13/carry[5] ), .IN2(n9), .Q(N1579) );
  OR2X1 U153 ( .IN1(a[27]), .IN2(\sub_114_I13/carry[4] ), .Q(
        \sub_114_I13/carry[5] ) );
  XNOR2X1 U154 ( .IN1(\sub_114_I13/carry[4] ), .IN2(a[27]), .Q(N1578) );
  AND2X1 U155 ( .IN1(N1116), .IN2(N2037), .Q(\sub_114_I13/carry[4] ) );
  XOR2X1 U156 ( .IN1(n3), .IN2(n20), .Q(N1577) );
  XNOR2X1 U157 ( .IN1(a[30]), .IN2(\sub_114_I11/carry[7] ), .Q(N1351) );
  OR2X1 U158 ( .IN1(n10), .IN2(\sub_114_I11/carry[6] ), .Q(
        \sub_114_I11/carry[7] ) );
  XNOR2X1 U159 ( .IN1(\sub_114_I11/carry[6] ), .IN2(n11), .Q(N1350) );
  OR2X1 U160 ( .IN1(n9), .IN2(\sub_114_I11/carry[5] ), .Q(
        \sub_114_I11/carry[6] ) );
  XNOR2X1 U161 ( .IN1(\sub_114_I11/carry[5] ), .IN2(n9), .Q(N1349) );
  OR2X1 U162 ( .IN1(a[27]), .IN2(\sub_114_I11/carry[4] ), .Q(
        \sub_114_I11/carry[5] ) );
  XNOR2X1 U163 ( .IN1(\sub_114_I11/carry[4] ), .IN2(a[27]), .Q(N1348) );
  AND2X1 U164 ( .IN1(\sub_114_I11/carry[3] ), .IN2(N2037), .Q(
        \sub_114_I11/carry[4] ) );
  XOR2X1 U165 ( .IN1(n2), .IN2(\sub_114_I11/carry[3] ), .Q(N1347) );
  OR2X1 U166 ( .IN1(N1116), .IN2(n5), .Q(\sub_114_I11/carry[3] ) );
  XNOR2X1 U167 ( .IN1(N662), .IN2(N1116), .Q(N1346) );
  XNOR2X1 U168 ( .IN1(a[30]), .IN2(\sub_114_I16/carry[7] ), .Q(N1926) );
  OR2X1 U169 ( .IN1(n10), .IN2(\sub_114_I16/carry[6] ), .Q(
        \sub_114_I16/carry[7] ) );
  XNOR2X1 U170 ( .IN1(\sub_114_I16/carry[6] ), .IN2(n11), .Q(N1925) );
  OR2X1 U171 ( .IN1(n9), .IN2(\sub_114_I16/carry[5] ), .Q(
        \sub_114_I16/carry[6] ) );
  XNOR2X1 U172 ( .IN1(\sub_114_I16/carry[5] ), .IN2(n9), .Q(N1924) );
  OR2X1 U173 ( .IN1(a[27]), .IN2(\sub_114_I16/carry[4] ), .Q(
        \sub_114_I16/carry[5] ) );
  XNOR2X1 U174 ( .IN1(\sub_114_I16/carry[4] ), .IN2(a[27]), .Q(N1923) );
  AND2X1 U175 ( .IN1(\sub_114_I16/carry[3] ), .IN2(n2), .Q(
        \sub_114_I16/carry[4] ) );
  XOR2X1 U176 ( .IN1(n3), .IN2(\sub_114_I16/carry[3] ), .Q(N1922) );
  AND2X1 U177 ( .IN1(\sub_114_I16/carry[2] ), .IN2(N1116), .Q(
        \sub_114_I16/carry[3] ) );
  XOR2X1 U178 ( .IN1(n20), .IN2(\sub_114_I16/carry[2] ), .Q(N1921) );
  AND2X1 U179 ( .IN1(N436), .IN2(N662), .Q(\sub_114_I16/carry[2] ) );
  XOR2X1 U180 ( .IN1(n4), .IN2(N436), .Q(N1920) );
  XNOR2X1 U181 ( .IN1(a[30]), .IN2(\sub_114_I10/carry[7] ), .Q(N1236) );
  OR2X1 U182 ( .IN1(n10), .IN2(\sub_114_I10/carry[6] ), .Q(
        \sub_114_I10/carry[7] ) );
  XNOR2X1 U183 ( .IN1(\sub_114_I10/carry[6] ), .IN2(n11), .Q(N1235) );
  OR2X1 U184 ( .IN1(n9), .IN2(\sub_114_I10/carry[5] ), .Q(
        \sub_114_I10/carry[6] ) );
  XNOR2X1 U185 ( .IN1(\sub_114_I10/carry[5] ), .IN2(n9), .Q(N1234) );
  OR2X1 U186 ( .IN1(n6), .IN2(\sub_114_I10/carry[4] ), .Q(
        \sub_114_I10/carry[5] ) );
  XNOR2X1 U187 ( .IN1(\sub_114_I10/carry[4] ), .IN2(n7), .Q(N1233) );
  AND2X1 U188 ( .IN1(\sub_114_I10/carry[3] ), .IN2(N2037), .Q(
        \sub_114_I10/carry[4] ) );
  XOR2X1 U189 ( .IN1(n2), .IN2(\sub_114_I10/carry[3] ), .Q(N1232) );
  OR2X1 U190 ( .IN1(N1116), .IN2(\sub_114_I10/carry[2] ), .Q(
        \sub_114_I10/carry[3] ) );
  XNOR2X1 U191 ( .IN1(\sub_114_I10/carry[2] ), .IN2(N1116), .Q(N1231) );
  OR2X1 U192 ( .IN1(N662), .IN2(N436), .Q(\sub_114_I10/carry[2] ) );
  XNOR2X1 U193 ( .IN1(N436), .IN2(n5), .Q(N1230) );
  XNOR2X1 U194 ( .IN1(a[30]), .IN2(\sub_114_I15/carry[7] ), .Q(N1811) );
  OR2X1 U195 ( .IN1(n10), .IN2(\sub_114_I15/carry[6] ), .Q(
        \sub_114_I15/carry[7] ) );
  XNOR2X1 U196 ( .IN1(\sub_114_I15/carry[6] ), .IN2(n10), .Q(N1810) );
  OR2X1 U197 ( .IN1(n9), .IN2(\sub_114_I15/carry[5] ), .Q(
        \sub_114_I15/carry[6] ) );
  XNOR2X1 U198 ( .IN1(\sub_114_I15/carry[5] ), .IN2(a[28]), .Q(N1809) );
  OR2X1 U199 ( .IN1(a[27]), .IN2(\sub_114_I15/carry[4] ), .Q(
        \sub_114_I15/carry[5] ) );
  XNOR2X1 U200 ( .IN1(\sub_114_I15/carry[4] ), .IN2(n7), .Q(N1808) );
  AND2X1 U201 ( .IN1(\sub_114_I15/carry[3] ), .IN2(N2037), .Q(
        \sub_114_I15/carry[4] ) );
  XOR2X1 U202 ( .IN1(n3), .IN2(\sub_114_I15/carry[3] ), .Q(N1807) );
  AND2X1 U203 ( .IN1(n4), .IN2(N1116), .Q(\sub_114_I15/carry[3] ) );
  XOR2X1 U204 ( .IN1(n20), .IN2(n5), .Q(N1806) );
  XNOR2X1 U205 ( .IN1(a[30]), .IN2(\sub_114_I14/carry[7] ), .Q(N1696) );
  OR2X1 U206 ( .IN1(n11), .IN2(\sub_114_I14/carry[6] ), .Q(
        \sub_114_I14/carry[7] ) );
  XNOR2X1 U207 ( .IN1(\sub_114_I14/carry[6] ), .IN2(n10), .Q(N1695) );
  OR2X1 U208 ( .IN1(n8), .IN2(\sub_114_I14/carry[5] ), .Q(
        \sub_114_I14/carry[6] ) );
  XNOR2X1 U209 ( .IN1(\sub_114_I14/carry[5] ), .IN2(n8), .Q(N1694) );
  OR2X1 U210 ( .IN1(n6), .IN2(\sub_114_I14/carry[4] ), .Q(
        \sub_114_I14/carry[5] ) );
  XNOR2X1 U211 ( .IN1(\sub_114_I14/carry[4] ), .IN2(n7), .Q(N1693) );
  AND2X1 U212 ( .IN1(\sub_114_I14/carry[3] ), .IN2(n2), .Q(
        \sub_114_I14/carry[4] ) );
  XOR2X1 U213 ( .IN1(n3), .IN2(\sub_114_I14/carry[3] ), .Q(N1692) );
  AND2X1 U214 ( .IN1(\sub_114_I14/carry[2] ), .IN2(N1116), .Q(
        \sub_114_I14/carry[3] ) );
  XOR2X1 U215 ( .IN1(n20), .IN2(\sub_114_I14/carry[2] ), .Q(N1691) );
  OR2X1 U216 ( .IN1(N662), .IN2(N436), .Q(\sub_114_I14/carry[2] ) );
  XNOR2X1 U217 ( .IN1(N436), .IN2(n5), .Q(N1690) );
  XNOR2X1 U218 ( .IN1(a[30]), .IN2(\sub_114_I8/carry[7] ), .Q(N1007) );
  OR2X1 U219 ( .IN1(n11), .IN2(\sub_114_I8/carry[6] ), .Q(
        \sub_114_I8/carry[7] ) );
  XNOR2X1 U220 ( .IN1(\sub_114_I8/carry[6] ), .IN2(n10), .Q(N1006) );
  OR2X1 U221 ( .IN1(n8), .IN2(\sub_114_I8/carry[5] ), .Q(\sub_114_I8/carry[6] ) );
  XNOR2X1 U222 ( .IN1(\sub_114_I8/carry[5] ), .IN2(a[28]), .Q(N1005) );
  OR2X1 U223 ( .IN1(n6), .IN2(\sub_114_I8/carry[4] ), .Q(\sub_114_I8/carry[5] ) );
  XNOR2X1 U224 ( .IN1(\sub_114_I8/carry[4] ), .IN2(n7), .Q(N1004) );
  OR2X1 U225 ( .IN1(N2037), .IN2(\sub_114_I8/carry[3] ), .Q(
        \sub_114_I8/carry[4] ) );
  XNOR2X1 U226 ( .IN1(\sub_114_I8/carry[3] ), .IN2(n3), .Q(N1003) );
  AND2X1 U227 ( .IN1(\sub_114_I8/carry[2] ), .IN2(N1116), .Q(
        \sub_114_I8/carry[3] ) );
  XOR2X1 U228 ( .IN1(n20), .IN2(\sub_114_I8/carry[2] ), .Q(N1002) );
  AND2X1 U229 ( .IN1(N436), .IN2(N662), .Q(\sub_114_I8/carry[2] ) );
  XOR2X1 U230 ( .IN1(n4), .IN2(N436), .Q(N1001) );
  XNOR2X1 U231 ( .IN1(a[30]), .IN2(\sub_114_I7/carry[7] ), .Q(N894) );
  OR2X1 U232 ( .IN1(n11), .IN2(\sub_114_I7/carry[6] ), .Q(
        \sub_114_I7/carry[7] ) );
  XNOR2X1 U233 ( .IN1(\sub_114_I7/carry[6] ), .IN2(n10), .Q(N893) );
  OR2X1 U234 ( .IN1(a[28]), .IN2(\sub_114_I7/carry[5] ), .Q(
        \sub_114_I7/carry[6] ) );
  XNOR2X1 U235 ( .IN1(\sub_114_I7/carry[5] ), .IN2(n8), .Q(N892) );
  OR2X1 U236 ( .IN1(n6), .IN2(\sub_114_I7/carry[4] ), .Q(\sub_114_I7/carry[5] ) );
  XNOR2X1 U237 ( .IN1(\sub_114_I7/carry[4] ), .IN2(n7), .Q(N891) );
  OR2X1 U238 ( .IN1(N2037), .IN2(\sub_114_I7/carry[3] ), .Q(
        \sub_114_I7/carry[4] ) );
  XNOR2X1 U239 ( .IN1(\sub_114_I7/carry[3] ), .IN2(n3), .Q(N890) );
  AND2X1 U240 ( .IN1(N662), .IN2(N1116), .Q(\sub_114_I7/carry[3] ) );
  XOR2X1 U241 ( .IN1(n20), .IN2(n5), .Q(N889) );
  XNOR2X1 U242 ( .IN1(a[30]), .IN2(\sub_114_I9/carry[7] ), .Q(N1121) );
  OR2X1 U243 ( .IN1(n11), .IN2(\sub_114_I9/carry[6] ), .Q(
        \sub_114_I9/carry[7] ) );
  XNOR2X1 U244 ( .IN1(\sub_114_I9/carry[6] ), .IN2(n10), .Q(N1120) );
  OR2X1 U245 ( .IN1(a[28]), .IN2(\sub_114_I9/carry[5] ), .Q(
        \sub_114_I9/carry[6] ) );
  XNOR2X1 U246 ( .IN1(\sub_114_I9/carry[5] ), .IN2(a[28]), .Q(N1119) );
  OR2X1 U247 ( .IN1(n6), .IN2(n2), .Q(\sub_114_I9/carry[5] ) );
  XNOR2X1 U248 ( .IN1(N2037), .IN2(n7), .Q(N1118) );
  XNOR2X1 U249 ( .IN1(a[30]), .IN2(\sub_114_I5/carry[7] ), .Q(N668) );
  OR2X1 U250 ( .IN1(n11), .IN2(\sub_114_I5/carry[6] ), .Q(
        \sub_114_I5/carry[7] ) );
  XNOR2X1 U251 ( .IN1(\sub_114_I5/carry[6] ), .IN2(n10), .Q(N667) );
  OR2X1 U252 ( .IN1(a[28]), .IN2(\sub_114_I5/carry[5] ), .Q(
        \sub_114_I5/carry[6] ) );
  XNOR2X1 U253 ( .IN1(\sub_114_I5/carry[5] ), .IN2(n8), .Q(N666) );
  OR2X1 U254 ( .IN1(n6), .IN2(\sub_114_I5/carry[4] ), .Q(\sub_114_I5/carry[5] ) );
  XNOR2X1 U255 ( .IN1(\sub_114_I5/carry[4] ), .IN2(n7), .Q(N665) );
  OR2X1 U256 ( .IN1(n2), .IN2(N1116), .Q(\sub_114_I5/carry[4] ) );
  XNOR2X1 U257 ( .IN1(N1116), .IN2(n3), .Q(N664) );
  XNOR2X1 U258 ( .IN1(a[30]), .IN2(\sub_114_I6/carry[7] ), .Q(N781) );
  OR2X1 U259 ( .IN1(n11), .IN2(\sub_114_I6/carry[6] ), .Q(
        \sub_114_I6/carry[7] ) );
  XNOR2X1 U260 ( .IN1(\sub_114_I6/carry[6] ), .IN2(n10), .Q(N780) );
  OR2X1 U261 ( .IN1(a[28]), .IN2(\sub_114_I6/carry[5] ), .Q(
        \sub_114_I6/carry[6] ) );
  XNOR2X1 U262 ( .IN1(\sub_114_I6/carry[5] ), .IN2(a[28]), .Q(N779) );
  OR2X1 U263 ( .IN1(a[27]), .IN2(\sub_114_I6/carry[4] ), .Q(
        \sub_114_I6/carry[5] ) );
  XNOR2X1 U264 ( .IN1(\sub_114_I6/carry[4] ), .IN2(n7), .Q(N778) );
  OR2X1 U265 ( .IN1(n2), .IN2(\sub_114_I6/carry[3] ), .Q(\sub_114_I6/carry[4] ) );
  XNOR2X1 U266 ( .IN1(\sub_114_I6/carry[3] ), .IN2(n3), .Q(N777) );
  AND2X1 U267 ( .IN1(\sub_114_I6/carry[2] ), .IN2(N1116), .Q(
        \sub_114_I6/carry[3] ) );
  XOR2X1 U268 ( .IN1(n20), .IN2(\sub_114_I6/carry[2] ), .Q(N776) );
  OR2X1 U269 ( .IN1(n4), .IN2(N436), .Q(\sub_114_I6/carry[2] ) );
  XNOR2X1 U270 ( .IN1(N436), .IN2(n5), .Q(N775) );
  XNOR2X1 U271 ( .IN1(a[30]), .IN2(\sub_114_I4/carry[7] ), .Q(N555) );
  OR2X1 U272 ( .IN1(a[29]), .IN2(\sub_114_I4/carry[6] ), .Q(
        \sub_114_I4/carry[7] ) );
  XNOR2X1 U273 ( .IN1(\sub_114_I4/carry[6] ), .IN2(n10), .Q(N554) );
  OR2X1 U274 ( .IN1(n8), .IN2(\sub_114_I4/carry[5] ), .Q(\sub_114_I4/carry[6] ) );
  XNOR2X1 U275 ( .IN1(\sub_114_I4/carry[5] ), .IN2(n8), .Q(N553) );
  OR2X1 U276 ( .IN1(n6), .IN2(\sub_114_I4/carry[4] ), .Q(\sub_114_I4/carry[5] ) );
  XNOR2X1 U277 ( .IN1(\sub_114_I4/carry[4] ), .IN2(n7), .Q(N552) );
  OR2X1 U278 ( .IN1(n2), .IN2(\sub_114_I4/carry[3] ), .Q(\sub_114_I4/carry[4] ) );
  XNOR2X1 U279 ( .IN1(\sub_114_I4/carry[3] ), .IN2(n3), .Q(N551) );
  OR2X1 U280 ( .IN1(N1116), .IN2(\sub_114_I4/carry[2] ), .Q(
        \sub_114_I4/carry[3] ) );
  XNOR2X1 U281 ( .IN1(\sub_114_I4/carry[2] ), .IN2(n20), .Q(N550) );
  AND2X1 U282 ( .IN1(N436), .IN2(n4), .Q(\sub_114_I4/carry[2] ) );
  XOR2X1 U283 ( .IN1(n5), .IN2(N436), .Q(N549) );
  XNOR2X1 U284 ( .IN1(a[30]), .IN2(\sub_114_I2_aco/carry[7] ), .Q(N375) );
  OR2X1 U285 ( .IN1(a[29]), .IN2(\sub_114_I2_aco/carry[6] ), .Q(
        \sub_114_I2_aco/carry[7] ) );
  XNOR2X1 U286 ( .IN1(\sub_114_I2_aco/carry[6] ), .IN2(n10), .Q(N374) );
  OR2X1 U287 ( .IN1(n8), .IN2(\sub_114_I2_aco/carry[5] ), .Q(
        \sub_114_I2_aco/carry[6] ) );
  XNOR2X1 U288 ( .IN1(\sub_114_I2_aco/carry[5] ), .IN2(a[28]), .Q(N373) );
  OR2X1 U289 ( .IN1(a[27]), .IN2(\sub_114_I2_aco/carry[4] ), .Q(
        \sub_114_I2_aco/carry[5] ) );
  XNOR2X1 U290 ( .IN1(\sub_114_I2_aco/carry[4] ), .IN2(n7), .Q(N372) );
  OR2X1 U291 ( .IN1(n2), .IN2(\sub_114_I2_aco/carry[3] ), .Q(
        \sub_114_I2_aco/carry[4] ) );
  XNOR2X1 U292 ( .IN1(\sub_114_I2_aco/carry[3] ), .IN2(n3), .Q(N371) );
  OR2X1 U293 ( .IN1(N1116), .IN2(\sub_114_I2_aco/carry[2] ), .Q(
        \sub_114_I2_aco/carry[3] ) );
  XNOR2X1 U294 ( .IN1(\sub_114_I2_aco/carry[2] ), .IN2(n20), .Q(N370) );
  OR2X1 U295 ( .IN1(N662), .IN2(\sub_114_I2_aco/carry[1] ), .Q(
        \sub_114_I2_aco/carry[2] ) );
  XNOR2X1 U296 ( .IN1(\sub_114_I2_aco/carry[1] ), .IN2(n5), .Q(N369) );
  OR2X1 U297 ( .IN1(N436), .IN2(n121), .Q(\sub_114_I2_aco/carry[1] ) );
  XNOR2X1 U298 ( .IN1(n121), .IN2(N436), .Q(N368) );
  XNOR2X1 U299 ( .IN1(a[30]), .IN2(\sub_114_I3/carry[7] ), .Q(N443) );
  OR2X1 U300 ( .IN1(a[29]), .IN2(\sub_114_I3/carry[6] ), .Q(
        \sub_114_I3/carry[7] ) );
  XNOR2X1 U301 ( .IN1(\sub_114_I3/carry[6] ), .IN2(n10), .Q(N442) );
  OR2X1 U302 ( .IN1(n8), .IN2(\sub_114_I3/carry[5] ), .Q(\sub_114_I3/carry[6] ) );
  XNOR2X1 U303 ( .IN1(\sub_114_I3/carry[5] ), .IN2(n8), .Q(N441) );
  OR2X1 U304 ( .IN1(a[27]), .IN2(\sub_114_I3/carry[4] ), .Q(
        \sub_114_I3/carry[5] ) );
  XNOR2X1 U305 ( .IN1(\sub_114_I3/carry[4] ), .IN2(n7), .Q(N440) );
  OR2X1 U306 ( .IN1(N2037), .IN2(\sub_114_I3/carry[3] ), .Q(
        \sub_114_I3/carry[4] ) );
  XNOR2X1 U307 ( .IN1(\sub_114_I3/carry[3] ), .IN2(n3), .Q(N439) );
  OR2X1 U308 ( .IN1(N1116), .IN2(n5), .Q(\sub_114_I3/carry[3] ) );
  XNOR2X1 U309 ( .IN1(n4), .IN2(n20), .Q(N438) );
  XNOR2X1 U310 ( .IN1(a[30]), .IN2(\sub_114_I12/carry[7] ), .Q(N1466) );
  OR2X1 U311 ( .IN1(a[29]), .IN2(\sub_114_I12/carry[6] ), .Q(
        \sub_114_I12/carry[7] ) );
  XNOR2X1 U312 ( .IN1(\sub_114_I12/carry[6] ), .IN2(n10), .Q(N1465) );
  OR2X1 U313 ( .IN1(n8), .IN2(\sub_114_I12/carry[5] ), .Q(
        \sub_114_I12/carry[6] ) );
  XNOR2X1 U314 ( .IN1(\sub_114_I12/carry[5] ), .IN2(a[28]), .Q(N1464) );
  OR2X1 U315 ( .IN1(n6), .IN2(\sub_114_I12/carry[4] ), .Q(
        \sub_114_I12/carry[5] ) );
  XNOR2X1 U316 ( .IN1(\sub_114_I12/carry[4] ), .IN2(a[27]), .Q(N1463) );
  AND2X1 U317 ( .IN1(\sub_114_I12/carry[3] ), .IN2(n2), .Q(
        \sub_114_I12/carry[4] ) );
  XOR2X1 U318 ( .IN1(n3), .IN2(\sub_114_I12/carry[3] ), .Q(N1462) );
  OR2X1 U319 ( .IN1(N1116), .IN2(\sub_114_I12/carry[2] ), .Q(
        \sub_114_I12/carry[3] ) );
  XNOR2X1 U320 ( .IN1(\sub_114_I12/carry[2] ), .IN2(n20), .Q(N1461) );
  AND2X1 U321 ( .IN1(N436), .IN2(N662), .Q(\sub_114_I12/carry[2] ) );
  XOR2X1 U322 ( .IN1(n5), .IN2(N436), .Q(N1460) );
  AND2X1 U323 ( .IN1(n61), .IN2(b_in[29]), .Q(n44) );
  NOR2X0 U324 ( .IN1(n55), .IN2(a_in[23]), .QN(n37) );
  AND2X1 U325 ( .IN1(n56), .IN2(n37), .Q(n38) );
  OA222X1 U326 ( .IN1(b_in[25]), .IN2(n57), .IN3(b_in[24]), .IN4(n38), .IN5(
        n37), .IN6(n56), .Q(n39) );
  AO221X1 U327 ( .IN1(b_in[25]), .IN2(n57), .IN3(b_in[26]), .IN4(n58), .IN5(
        n39), .Q(n40) );
  OA221X1 U328 ( .IN1(b_in[27]), .IN2(n59), .IN3(b_in[26]), .IN4(n58), .IN5(
        n40), .Q(n41) );
  AO221X1 U329 ( .IN1(b_in[27]), .IN2(n59), .IN3(b_in[28]), .IN4(n60), .IN5(
        n41), .Q(n42) );
  OA221X1 U330 ( .IN1(b_in[29]), .IN2(n61), .IN3(b_in[28]), .IN4(n60), .IN5(
        n42), .Q(n43) );
  OA22X1 U331 ( .IN1(b_in[30]), .IN2(n62), .IN3(n44), .IN4(n43), .Q(n45) );
  AO21X1 U332 ( .IN1(b_in[30]), .IN2(n62), .IN3(n45), .Q(N54) );
  NOR2X0 U333 ( .IN1(n63), .IN2(n64), .QN(sum_31) );
  MUX21X1 U334 ( .IN1(n25), .IN2(n31), .S(N59), .Q(n64) );
  AO22X1 U335 ( .IN1(n12), .IN2(n66), .IN3(n67), .IN4(n68), .Q(sum[9]) );
  NOR2X0 U336 ( .IN1(n69), .IN2(n70), .QN(n67) );
  AO21X1 U337 ( .IN1(n65), .IN2(n71), .IN3(n72), .Q(sum[8]) );
  AND4X1 U338 ( .IN1(n73), .IN2(n74), .IN3(n75), .IN4(n76), .Q(n72) );
  AO22X1 U339 ( .IN1(n12), .IN2(n77), .IN3(n78), .IN4(n68), .Q(sum[7]) );
  NOR2X0 U340 ( .IN1(n79), .IN2(n80), .QN(n78) );
  NOR2X0 U341 ( .IN1(n84), .IN2(n85), .QN(n68) );
  AO21X1 U342 ( .IN1(n65), .IN2(n87), .IN3(n88), .Q(sum[5]) );
  NOR4X0 U343 ( .IN1(n89), .IN2(n90), .IN3(n91), .IN4(n84), .QN(n88) );
  AO22X1 U344 ( .IN1(n65), .IN2(n92), .IN3(n93), .IN4(n76), .Q(sum[4]) );
  NOR2X0 U345 ( .IN1(n94), .IN2(n95), .QN(n93) );
  AO21X1 U346 ( .IN1(n65), .IN2(n96), .IN3(n97), .Q(sum[3]) );
  NOR4X0 U347 ( .IN1(n98), .IN2(n99), .IN3(n100), .IN4(n84), .QN(n97) );
  AO22X1 U348 ( .IN1(n65), .IN2(n101), .IN3(n102), .IN4(n76), .Q(sum[2]) );
  NOR2X0 U349 ( .IN1(n103), .IN2(n104), .QN(n102) );
  NAND4X0 U350 ( .IN1(n76), .IN2(n105), .IN3(n106), .IN4(n107), .QN(sum[22])
         );
  NOR3X0 U351 ( .IN1(n95), .IN2(n108), .IN3(n109), .QN(n107) );
  AO22X1 U352 ( .IN1(n65), .IN2(n109), .IN3(n76), .IN4(n110), .Q(sum[21]) );
  NAND4X0 U353 ( .IN1(n111), .IN2(n112), .IN3(n113), .IN4(n114), .QN(n110) );
  NOR4X0 U354 ( .IN1(n115), .IN2(n116), .IN3(n117), .IN4(n118), .QN(n114) );
  MUX21X1 U355 ( .IN1(n119), .IN2(n120), .S(n121), .Q(n118) );
  NOR2X0 U356 ( .IN1(n122), .IN2(n123), .QN(n117) );
  AO222X1 U357 ( .IN1(n124), .IN2(n125), .IN3(n126), .IN4(n127), .IN5(n99), 
        .IN6(n128), .Q(n116) );
  AO221X1 U358 ( .IN1(n129), .IN2(n130), .IN3(n131), .IN4(n132), .IN5(n133), 
        .Q(n115) );
  AO222X1 U359 ( .IN1(n134), .IN2(n135), .IN3(n89), .IN4(n136), .IN5(n137), 
        .IN6(n138), .Q(n133) );
  INVX0 U360 ( .INP(n139), .ZN(n130) );
  OA221X1 U361 ( .IN1(n100), .IN2(n140), .IN3(n141), .IN4(n142), .IN5(n143), 
        .Q(n113) );
  OA222X1 U362 ( .IN1(n144), .IN2(n145), .IN3(n146), .IN4(n147), .IN5(n148), 
        .IN6(n149), .Q(n143) );
  INVX0 U363 ( .INP(n150), .ZN(n144) );
  OA222X1 U364 ( .IN1(n69), .IN2(n151), .IN3(n94), .IN4(n152), .IN5(n79), 
        .IN6(n73), .Q(n112) );
  OA222X1 U365 ( .IN1(n153), .IN2(n154), .IN3(n155), .IN4(n156), .IN5(n157), 
        .IN6(n158), .Q(n111) );
  AO22X1 U366 ( .IN1(n65), .IN2(n120), .IN3(n76), .IN4(n159), .Q(sum[20]) );
  NAND4X0 U367 ( .IN1(n160), .IN2(n161), .IN3(n162), .IN4(n163), .QN(n159) );
  NOR2X0 U368 ( .IN1(n164), .IN2(n165), .QN(n163) );
  OAI222X1 U369 ( .IN1(n166), .IN2(n167), .IN3(n154), .IN4(n168), .IN5(n149), 
        .IN6(n169), .QN(n165) );
  AO222X1 U370 ( .IN1(n170), .IN2(n81), .IN3(n90), .IN4(n171), .IN5(n134), 
        .IN6(n172), .Q(n164) );
  OA221X1 U371 ( .IN1(n79), .IN2(n156), .IN3(n122), .IN4(n173), .IN5(n174), 
        .Q(n162) );
  AOI222X1 U372 ( .IN1(n119), .IN2(n175), .IN3(n176), .IN4(n14), .IN5(n150), 
        .IN6(\sub_114_I2_aco/B[0] ), .QN(n174) );
  OA221X1 U373 ( .IN1(n148), .IN2(n178), .IN3(n153), .IN4(n179), .IN5(n180), 
        .Q(n161) );
  OA222X1 U374 ( .IN1(n181), .IN2(n182), .IN3(n183), .IN4(n147), .IN5(n184), 
        .IN6(n185), .Q(n180) );
  INVX0 U375 ( .INP(n186), .ZN(n153) );
  INVX0 U376 ( .INP(n187), .ZN(n148) );
  OA221X1 U377 ( .IN1(n94), .IN2(n83), .IN3(n188), .IN4(n123), .IN5(n189), .Q(
        n160) );
  OA222X1 U378 ( .IN1(n190), .IN2(n140), .IN3(n155), .IN4(n151), .IN5(n191), 
        .IN6(n158), .Q(n189) );
  INVX0 U379 ( .INP(n192), .ZN(n94) );
  AO21X1 U380 ( .IN1(n65), .IN2(n193), .IN3(n194), .Q(sum[1]) );
  NOR4X0 U381 ( .IN1(n108), .IN2(n104), .IN3(n122), .IN4(n84), .QN(n194) );
  INVX0 U382 ( .INP(n105), .ZN(n104) );
  AO22X1 U383 ( .IN1(n65), .IN2(n119), .IN3(n76), .IN4(n195), .Q(sum[19]) );
  NAND4X0 U384 ( .IN1(n196), .IN2(n197), .IN3(n198), .IN4(n199), .QN(n195) );
  OA221X1 U385 ( .IN1(n200), .IN2(n149), .IN3(n201), .IN4(n151), .IN5(n202), 
        .Q(n199) );
  OA222X1 U386 ( .IN1(n191), .IN2(n73), .IN3(n190), .IN4(n152), .IN5(n203), 
        .IN6(n158), .Q(n202) );
  OA221X1 U387 ( .IN1(n157), .IN2(n156), .IN3(n204), .IN4(n205), .IN5(n206), 
        .Q(n198) );
  OA22X1 U388 ( .IN1(n147), .IN2(n69), .IN3(n207), .IN4(n185), .Q(n206) );
  INVX0 U389 ( .INP(n208), .ZN(n204) );
  OA221X1 U390 ( .IN1(n209), .IN2(n166), .IN3(n210), .IN4(n182), .IN5(n211), 
        .Q(n197) );
  OA22X1 U391 ( .IN1(n212), .IN2(n154), .IN3(n168), .IN4(n179), .Q(n211) );
  OA221X1 U392 ( .IN1(n213), .IN2(n140), .IN3(n188), .IN4(n173), .IN5(n214), 
        .Q(n196) );
  OA21X1 U393 ( .IN1(n215), .IN2(n83), .IN3(n216), .Q(n214) );
  MUX21X1 U394 ( .IN1(n169), .IN2(n217), .S(n178), .Q(n216) );
  INVX0 U395 ( .INP(n218), .ZN(n217) );
  INVX0 U396 ( .INP(n219), .ZN(n169) );
  AO22X1 U397 ( .IN1(n65), .IN2(n150), .IN3(n76), .IN4(n220), .Q(sum[18]) );
  NAND4X0 U398 ( .IN1(n221), .IN2(n222), .IN3(n223), .IN4(n224), .QN(n220) );
  OA221X1 U399 ( .IN1(n201), .IN2(n205), .IN3(n215), .IN4(n158), .IN5(n225), 
        .Q(n224) );
  OA222X1 U400 ( .IN1(n226), .IN2(n151), .IN3(n203), .IN4(n73), .IN5(n213), 
        .IN6(n152), .Q(n225) );
  OA221X1 U401 ( .IN1(n227), .IN2(n147), .IN3(n191), .IN4(n156), .IN5(n228), 
        .Q(n223) );
  OA22X1 U402 ( .IN1(n229), .IN2(n154), .IN3(n200), .IN4(n178), .Q(n228) );
  INVX0 U403 ( .INP(n230), .ZN(n200) );
  OA221X1 U404 ( .IN1(n231), .IN2(n179), .IN3(n232), .IN4(n166), .IN5(n233), 
        .Q(n222) );
  AOI22X1 U405 ( .IN1(n234), .IN2(n235), .IN3(n125), .IN4(n236), .QN(n233) );
  OA221X1 U406 ( .IN1(n188), .IN2(n140), .IN3(n190), .IN4(n83), .IN5(n237), 
        .Q(n221) );
  OA22X1 U407 ( .IN1(n238), .IN2(n185), .IN3(n239), .IN4(n182), .Q(n237) );
  INVX0 U408 ( .INP(n240), .ZN(n190) );
  NAND4X0 U409 ( .IN1(n242), .IN2(n243), .IN3(n244), .IN4(n245), .QN(n241) );
  OA221X1 U410 ( .IN1(n213), .IN2(n83), .IN3(n188), .IN4(n152), .IN5(n246), 
        .Q(n245) );
  OA22X1 U411 ( .IN1(n247), .IN2(n158), .IN3(n203), .IN4(n156), .Q(n246) );
  INVX0 U412 ( .INP(n248), .ZN(n213) );
  OA222X1 U413 ( .IN1(n249), .IN2(n154), .IN3(n226), .IN4(n205), .IN5(n147), 
        .IN6(n201), .Q(n244) );
  OA222X1 U414 ( .IN1(n238), .IN2(n182), .IN3(n227), .IN4(n185), .IN5(n215), 
        .IN6(n73), .Q(n243) );
  OA221X1 U415 ( .IN1(n191), .IN2(n151), .IN3(n250), .IN4(n166), .IN5(n251), 
        .Q(n242) );
  INVX0 U416 ( .INP(n252), .ZN(n251) );
  MUX21X1 U417 ( .IN1(n253), .IN2(n254), .S(n179), .Q(n252) );
  INVX0 U418 ( .INP(n255), .ZN(n191) );
  AO22X1 U419 ( .IN1(n12), .IN2(n256), .IN3(n76), .IN4(n257), .Q(sum[16]) );
  NAND4X0 U420 ( .IN1(n258), .IN2(n259), .IN3(n260), .IN4(n261), .QN(n257) );
  OA221X1 U421 ( .IN1(n188), .IN2(n83), .IN3(n262), .IN4(n158), .IN5(n263), 
        .Q(n261) );
  OA22X1 U422 ( .IN1(n247), .IN2(n73), .IN3(n264), .IN4(n156), .Q(n263) );
  INVX0 U423 ( .INP(n265), .ZN(n188) );
  OA222X1 U424 ( .IN1(n249), .IN2(n179), .IN3(n203), .IN4(n151), .IN5(n185), 
        .IN6(n201), .Q(n260) );
  INVX0 U425 ( .INP(n266), .ZN(n201) );
  AOI222X1 U426 ( .IN1(n127), .IN2(n267), .IN3(n268), .IN4(n134), .IN5(n269), 
        .IN6(n270), .QN(n259) );
  INVX0 U427 ( .INP(n271), .ZN(n268) );
  OA222X1 U428 ( .IN1(n147), .IN2(n226), .IN3(n272), .IN4(n182), .IN5(n273), 
        .IN6(n166), .Q(n258) );
  INVX0 U429 ( .INP(n274), .ZN(n226) );
  AO22X1 U430 ( .IN1(n12), .IN2(n275), .IN3(n76), .IN4(n276), .Q(sum[15]) );
  NAND4X0 U431 ( .IN1(n277), .IN2(n278), .IN3(n279), .IN4(n280), .QN(n276) );
  OA221X1 U432 ( .IN1(n281), .IN2(n158), .IN3(n264), .IN4(n151), .IN5(n282), 
        .Q(n280) );
  OA222X1 U433 ( .IN1(n283), .IN2(n185), .IN3(n247), .IN4(n156), .IN5(n262), 
        .IN6(n73), .Q(n282) );
  OA22X1 U434 ( .IN1(n147), .IN2(n271), .IN3(n203), .IN4(n205), .Q(n279) );
  OR2X1 U435 ( .IN1(n182), .IN2(n284), .Q(n278) );
  MUX21X1 U436 ( .IN1(n285), .IN2(n286), .S(n166), .Q(n277) );
  INVX0 U437 ( .INP(n287), .ZN(n286) );
  AO22X1 U438 ( .IN1(n12), .IN2(n288), .IN3(n76), .IN4(n289), .Q(sum[14]) );
  NAND4X0 U439 ( .IN1(n290), .IN2(n291), .IN3(n292), .IN4(n293), .QN(n289) );
  OA222X1 U440 ( .IN1(n262), .IN2(n156), .IN3(n247), .IN4(n151), .IN5(n264), 
        .IN6(n205), .Q(n293) );
  OA22X1 U441 ( .IN1(n283), .IN2(n182), .IN3(n294), .IN4(n295), .Q(n292) );
  OA22X1 U442 ( .IN1(n147), .IN2(n203), .IN3(n296), .IN4(n166), .Q(n291) );
  OA22X1 U443 ( .IN1(n281), .IN2(n73), .IN3(n185), .IN4(n271), .Q(n290) );
  AO22X1 U444 ( .IN1(n12), .IN2(n297), .IN3(n76), .IN4(n298), .Q(sum[13]) );
  NAND3X0 U445 ( .IN1(n299), .IN2(n300), .IN3(n301), .QN(n298) );
  OA222X1 U446 ( .IN1(n262), .IN2(n151), .IN3(n302), .IN4(n156), .IN5(n247), 
        .IN6(n205), .Q(n301) );
  NAND2X0 U447 ( .IN1(n303), .IN2(n304), .QN(n300) );
  MUX21X1 U448 ( .IN1(n203), .IN2(n305), .S(n185), .Q(n299) );
  AO22X1 U449 ( .IN1(n12), .IN2(n306), .IN3(n76), .IN4(n307), .Q(sum[12]) );
  AO221X1 U450 ( .IN1(n134), .IN2(n308), .IN3(n309), .IN4(n310), .IN5(n311), 
        .Q(n307) );
  MUX21X1 U451 ( .IN1(n312), .IN2(n313), .S(n147), .Q(n311) );
  INVX0 U452 ( .INP(n247), .ZN(n312) );
  AO22X1 U453 ( .IN1(n12), .IN2(n314), .IN3(n76), .IN4(n315), .Q(sum[11]) );
  MUX21X1 U454 ( .IN1(n310), .IN2(n316), .S(n205), .Q(n315) );
  AO21X1 U455 ( .IN1(n65), .IN2(n317), .IN3(n318), .Q(sum[10]) );
  NOR4X0 U456 ( .IN1(n134), .IN2(n309), .IN3(n84), .IN4(n319), .QN(n318) );
  AO22X1 U457 ( .IN1(n12), .IN2(n320), .IN3(n321), .IN4(n76), .Q(sum[0]) );
  INVX0 U458 ( .INP(n84), .ZN(n76) );
  AO21X1 U459 ( .IN1(n322), .IN2(n323), .IN3(n65), .Q(n84) );
  NOR2X0 U460 ( .IN1(n108), .IN2(n141), .QN(n321) );
  INVX0 U461 ( .INP(n142), .ZN(n108) );
  MUX21X1 U462 ( .IN1(b_in[9]), .IN2(a_in[9]), .S(n32), .Q(b[9]) );
  MUX21X1 U463 ( .IN1(b_in[8]), .IN2(a_in[8]), .S(n32), .Q(b[8]) );
  MUX21X1 U464 ( .IN1(b_in[7]), .IN2(a_in[7]), .S(n32), .Q(b[7]) );
  MUX21X1 U465 ( .IN1(b_in[6]), .IN2(a_in[6]), .S(n32), .Q(b[6]) );
  MUX21X1 U466 ( .IN1(b_in[5]), .IN2(a_in[5]), .S(n32), .Q(b[5]) );
  MUX21X1 U467 ( .IN1(b_in[4]), .IN2(a_in[4]), .S(n32), .Q(b[4]) );
  MUX21X1 U468 ( .IN1(b_in[3]), .IN2(a_in[3]), .S(n32), .Q(b[3]) );
  MUX21X1 U469 ( .IN1(b_in[30]), .IN2(a_in[30]), .S(n32), .Q(b[30]) );
  MUX21X1 U470 ( .IN1(b_in[2]), .IN2(a_in[2]), .S(n32), .Q(b[2]) );
  MUX21X1 U471 ( .IN1(b_in[29]), .IN2(a_in[29]), .S(n32), .Q(b[29]) );
  MUX21X1 U472 ( .IN1(b_in[28]), .IN2(a_in[28]), .S(n32), .Q(b[28]) );
  MUX21X1 U473 ( .IN1(b_in[27]), .IN2(a_in[27]), .S(n32), .Q(b[27]) );
  MUX21X1 U474 ( .IN1(b_in[26]), .IN2(a_in[26]), .S(n33), .Q(b[26]) );
  MUX21X1 U475 ( .IN1(b_in[25]), .IN2(a_in[25]), .S(n33), .Q(b[25]) );
  MUX21X1 U476 ( .IN1(b_in[24]), .IN2(a_in[24]), .S(n33), .Q(b[24]) );
  MUX21X1 U477 ( .IN1(b_in[23]), .IN2(a_in[23]), .S(n33), .Q(b[23]) );
  MUX21X1 U478 ( .IN1(b_in[22]), .IN2(a_in[22]), .S(n33), .Q(b[22]) );
  MUX21X1 U479 ( .IN1(b_in[21]), .IN2(a_in[21]), .S(n33), .Q(b[21]) );
  MUX21X1 U480 ( .IN1(b_in[20]), .IN2(a_in[20]), .S(n33), .Q(b[20]) );
  MUX21X1 U481 ( .IN1(b_in[1]), .IN2(a_in[1]), .S(n33), .Q(b[1]) );
  MUX21X1 U482 ( .IN1(b_in[19]), .IN2(a_in[19]), .S(n33), .Q(b[19]) );
  MUX21X1 U483 ( .IN1(b_in[18]), .IN2(a_in[18]), .S(n33), .Q(b[18]) );
  MUX21X1 U484 ( .IN1(b_in[17]), .IN2(a_in[17]), .S(n33), .Q(b[17]) );
  MUX21X1 U485 ( .IN1(b_in[16]), .IN2(a_in[16]), .S(n33), .Q(b[16]) );
  MUX21X1 U486 ( .IN1(b_in[15]), .IN2(a_in[15]), .S(n34), .Q(b[15]) );
  MUX21X1 U487 ( .IN1(b_in[14]), .IN2(a_in[14]), .S(n34), .Q(b[14]) );
  MUX21X1 U488 ( .IN1(b_in[13]), .IN2(a_in[13]), .S(n34), .Q(b[13]) );
  MUX21X1 U489 ( .IN1(b_in[12]), .IN2(a_in[12]), .S(n34), .Q(b[12]) );
  MUX21X1 U490 ( .IN1(b_in[11]), .IN2(a_in[11]), .S(n34), .Q(b[11]) );
  MUX21X1 U491 ( .IN1(b_in[10]), .IN2(a_in[10]), .S(n34), .Q(b[10]) );
  MUX21X1 U492 ( .IN1(b_in[0]), .IN2(a_in[0]), .S(n34), .Q(b[0]) );
  MUX21X1 U493 ( .IN1(a_in[9]), .IN2(b_in[9]), .S(n34), .Q(a[9]) );
  MUX21X1 U494 ( .IN1(a_in[8]), .IN2(b_in[8]), .S(n34), .Q(a[8]) );
  MUX21X1 U495 ( .IN1(a_in[7]), .IN2(b_in[7]), .S(n34), .Q(a[7]) );
  MUX21X1 U496 ( .IN1(a_in[6]), .IN2(b_in[6]), .S(n34), .Q(a[6]) );
  MUX21X1 U497 ( .IN1(a_in[5]), .IN2(b_in[5]), .S(n34), .Q(a[5]) );
  MUX21X1 U498 ( .IN1(a_in[4]), .IN2(b_in[4]), .S(n35), .Q(a[4]) );
  MUX21X1 U499 ( .IN1(a_in[3]), .IN2(b_in[3]), .S(n35), .Q(a[3]) );
  MUX21X1 U500 ( .IN1(a_in[2]), .IN2(b_in[2]), .S(n35), .Q(a[2]) );
  MUX21X1 U501 ( .IN1(a_in[22]), .IN2(b_in[22]), .S(n35), .Q(a[22]) );
  MUX21X1 U502 ( .IN1(a_in[21]), .IN2(b_in[21]), .S(n35), .Q(a[21]) );
  MUX21X1 U503 ( .IN1(a_in[20]), .IN2(b_in[20]), .S(n35), .Q(a[20]) );
  MUX21X1 U504 ( .IN1(a_in[1]), .IN2(b_in[1]), .S(n35), .Q(a[1]) );
  MUX21X1 U505 ( .IN1(a_in[19]), .IN2(b_in[19]), .S(n35), .Q(a[19]) );
  MUX21X1 U506 ( .IN1(a_in[18]), .IN2(b_in[18]), .S(n35), .Q(a[18]) );
  MUX21X1 U507 ( .IN1(a_in[17]), .IN2(b_in[17]), .S(n35), .Q(a[17]) );
  MUX21X1 U508 ( .IN1(a_in[16]), .IN2(b_in[16]), .S(n35), .Q(a[16]) );
  MUX21X1 U509 ( .IN1(a_in[15]), .IN2(b_in[15]), .S(n35), .Q(a[15]) );
  MUX21X1 U510 ( .IN1(a_in[14]), .IN2(b_in[14]), .S(N54), .Q(a[14]) );
  MUX21X1 U511 ( .IN1(a_in[13]), .IN2(b_in[13]), .S(n36), .Q(a[13]) );
  MUX21X1 U512 ( .IN1(a_in[12]), .IN2(b_in[12]), .S(N54), .Q(a[12]) );
  MUX21X1 U513 ( .IN1(a_in[11]), .IN2(b_in[11]), .S(n36), .Q(a[11]) );
  MUX21X1 U514 ( .IN1(a_in[10]), .IN2(b_in[10]), .S(N54), .Q(a[10]) );
  MUX21X1 U515 ( .IN1(a_in[0]), .IN2(b_in[0]), .S(n36), .Q(a[0]) );
  OR4X1 U516 ( .IN1(n325), .IN2(n326), .IN3(n327), .IN4(n328), .Q(N2810) );
  AO221X1 U517 ( .IN1(N2271), .IN2(n329), .IN3(N2616), .IN4(n330), .IN5(n331), 
        .Q(n328) );
  AO22X1 U518 ( .IN1(N297), .IN2(n12), .IN3(N2731), .IN4(n332), .Q(n331) );
  AO222X1 U519 ( .IN1(N2156), .IN2(n333), .IN3(N2501), .IN4(n334), .IN5(N2041), 
        .IN6(n335), .Q(n327) );
  AND2X1 U520 ( .IN1(N2386), .IN2(n336), .Q(n326) );
  OA21X1 U521 ( .IN1(n337), .IN2(n338), .IN3(n339), .Q(n325) );
  AO221X1 U522 ( .IN1(N1236), .IN2(n137), .IN3(N1926), .IN4(n340), .IN5(n341), 
        .Q(n338) );
  AO22X1 U523 ( .IN1(N1351), .IN2(n304), .IN3(N1581), .IN4(n309), .Q(n341) );
  AO221X1 U524 ( .IN1(N1466), .IN2(n134), .IN3(n342), .IN4(n343), .IN5(n344), 
        .Q(n337) );
  AO22X1 U525 ( .IN1(N1696), .IN2(n85), .IN3(N1811), .IN4(n170), .Q(n344) );
  OR2X1 U526 ( .IN1(n345), .IN2(n346), .Q(n343) );
  AO221X1 U527 ( .IN1(N668), .IN2(n235), .IN3(N1121), .IN4(n129), .IN5(n347), 
        .Q(n346) );
  AO22X1 U528 ( .IN1(N894), .IN2(n270), .IN3(N1007), .IN4(n131), .Q(n347) );
  AO221X1 U529 ( .IN1(N443), .IN2(n14), .IN3(N375), .IN4(n348), .IN5(n349), 
        .Q(n345) );
  AO22X1 U530 ( .IN1(N555), .IN2(n124), .IN3(N781), .IN4(n126), .Q(n349) );
  OR4X1 U531 ( .IN1(n350), .IN2(n351), .IN3(n352), .IN4(n353), .Q(N2809) );
  AO221X1 U532 ( .IN1(N2270), .IN2(n329), .IN3(N2615), .IN4(n330), .IN5(n354), 
        .Q(n353) );
  AO22X1 U533 ( .IN1(N296), .IN2(n12), .IN3(N2730), .IN4(n332), .Q(n354) );
  AO222X1 U534 ( .IN1(N2155), .IN2(n333), .IN3(N2500), .IN4(n334), .IN5(N2040), 
        .IN6(n335), .Q(n352) );
  AND2X1 U535 ( .IN1(N2385), .IN2(n336), .Q(n351) );
  OA21X1 U536 ( .IN1(n355), .IN2(n356), .IN3(n339), .Q(n350) );
  AO221X1 U537 ( .IN1(N1235), .IN2(n137), .IN3(N1925), .IN4(n340), .IN5(n357), 
        .Q(n356) );
  AO22X1 U538 ( .IN1(N1350), .IN2(n304), .IN3(N1580), .IN4(n309), .Q(n357) );
  AO221X1 U539 ( .IN1(N1465), .IN2(n134), .IN3(n342), .IN4(n358), .IN5(n359), 
        .Q(n355) );
  AO22X1 U540 ( .IN1(N1695), .IN2(n85), .IN3(N1810), .IN4(n170), .Q(n359) );
  OR2X1 U541 ( .IN1(n360), .IN2(n361), .Q(n358) );
  AO221X1 U542 ( .IN1(N667), .IN2(n235), .IN3(N1120), .IN4(n129), .IN5(n362), 
        .Q(n361) );
  AO22X1 U543 ( .IN1(N893), .IN2(n270), .IN3(N1006), .IN4(n131), .Q(n362) );
  AO221X1 U544 ( .IN1(N442), .IN2(n14), .IN3(N374), .IN4(n348), .IN5(n363), 
        .Q(n360) );
  AO22X1 U545 ( .IN1(N554), .IN2(n124), .IN3(N780), .IN4(n126), .Q(n363) );
  OR4X1 U546 ( .IN1(n364), .IN2(n365), .IN3(n366), .IN4(n367), .Q(N2808) );
  AO221X1 U547 ( .IN1(N2269), .IN2(n329), .IN3(N2614), .IN4(n330), .IN5(n368), 
        .Q(n367) );
  AO22X1 U548 ( .IN1(N295), .IN2(n12), .IN3(N2729), .IN4(n332), .Q(n368) );
  AO222X1 U549 ( .IN1(N2154), .IN2(n333), .IN3(N2499), .IN4(n334), .IN5(N2039), 
        .IN6(n335), .Q(n366) );
  AND2X1 U550 ( .IN1(N2384), .IN2(n336), .Q(n365) );
  OA21X1 U551 ( .IN1(n369), .IN2(n370), .IN3(n339), .Q(n364) );
  AO221X1 U552 ( .IN1(N1234), .IN2(n137), .IN3(N1924), .IN4(n340), .IN5(n371), 
        .Q(n370) );
  AO22X1 U553 ( .IN1(N1349), .IN2(n304), .IN3(N1579), .IN4(n309), .Q(n371) );
  AO221X1 U554 ( .IN1(N1464), .IN2(n134), .IN3(n342), .IN4(n372), .IN5(n373), 
        .Q(n369) );
  AO22X1 U555 ( .IN1(N1694), .IN2(n85), .IN3(N1809), .IN4(n170), .Q(n373) );
  OR2X1 U556 ( .IN1(n374), .IN2(n375), .Q(n372) );
  AO221X1 U557 ( .IN1(N666), .IN2(n235), .IN3(N1119), .IN4(n129), .IN5(n376), 
        .Q(n375) );
  AO22X1 U558 ( .IN1(N892), .IN2(n270), .IN3(N1005), .IN4(n131), .Q(n376) );
  AO221X1 U559 ( .IN1(N441), .IN2(n14), .IN3(N373), .IN4(n348), .IN5(n377), 
        .Q(n374) );
  AO22X1 U560 ( .IN1(N553), .IN2(n124), .IN3(N779), .IN4(n126), .Q(n377) );
  OR4X1 U561 ( .IN1(n378), .IN2(n379), .IN3(n380), .IN4(n381), .Q(N2807) );
  AO221X1 U562 ( .IN1(N2268), .IN2(n329), .IN3(N2613), .IN4(n330), .IN5(n382), 
        .Q(n381) );
  AO22X1 U563 ( .IN1(N294), .IN2(n12), .IN3(N2728), .IN4(n332), .Q(n382) );
  AO222X1 U564 ( .IN1(N2153), .IN2(n333), .IN3(N2498), .IN4(n334), .IN5(n26), 
        .IN6(n335), .Q(n380) );
  AND2X1 U565 ( .IN1(N2383), .IN2(n336), .Q(n379) );
  OA21X1 U566 ( .IN1(n383), .IN2(n384), .IN3(n339), .Q(n378) );
  AO221X1 U567 ( .IN1(N1233), .IN2(n137), .IN3(N1923), .IN4(n340), .IN5(n385), 
        .Q(n384) );
  AO22X1 U568 ( .IN1(N1348), .IN2(n304), .IN3(N1578), .IN4(n309), .Q(n385) );
  AO221X1 U569 ( .IN1(N1463), .IN2(n134), .IN3(n342), .IN4(n386), .IN5(n387), 
        .Q(n383) );
  AO22X1 U570 ( .IN1(N1693), .IN2(n85), .IN3(N1808), .IN4(n170), .Q(n387) );
  OR2X1 U571 ( .IN1(n388), .IN2(n389), .Q(n386) );
  AO221X1 U572 ( .IN1(N665), .IN2(n235), .IN3(N1118), .IN4(n129), .IN5(n390), 
        .Q(n389) );
  AO22X1 U573 ( .IN1(N891), .IN2(n270), .IN3(N1004), .IN4(n131), .Q(n390) );
  AO22X1 U574 ( .IN1(N552), .IN2(n124), .IN3(N778), .IN4(n126), .Q(n391) );
  OR4X1 U575 ( .IN1(n392), .IN2(n393), .IN3(n394), .IN4(n395), .Q(N2806) );
  AO221X1 U576 ( .IN1(N2267), .IN2(n329), .IN3(N2612), .IN4(n330), .IN5(n396), 
        .Q(n395) );
  AO22X1 U577 ( .IN1(N293), .IN2(n12), .IN3(N2727), .IN4(n332), .Q(n396) );
  AO222X1 U578 ( .IN1(N2152), .IN2(n333), .IN3(N2497), .IN4(n334), .IN5(n2), 
        .IN6(n335), .Q(n394) );
  AND2X1 U579 ( .IN1(N2382), .IN2(n336), .Q(n393) );
  OA21X1 U580 ( .IN1(n397), .IN2(n398), .IN3(n339), .Q(n392) );
  AO221X1 U581 ( .IN1(N1232), .IN2(n137), .IN3(N1922), .IN4(n340), .IN5(n399), 
        .Q(n398) );
  AO22X1 U582 ( .IN1(N1347), .IN2(n304), .IN3(N1577), .IN4(n309), .Q(n399) );
  AO221X1 U583 ( .IN1(N1462), .IN2(n134), .IN3(n342), .IN4(n400), .IN5(n401), 
        .Q(n397) );
  AO22X1 U584 ( .IN1(N1692), .IN2(n85), .IN3(N1807), .IN4(n170), .Q(n401) );
  OR2X1 U585 ( .IN1(n402), .IN2(n403), .Q(n400) );
  AO221X1 U586 ( .IN1(N664), .IN2(n235), .IN3(n19), .IN4(n129), .IN5(n404), 
        .Q(n403) );
  AO22X1 U587 ( .IN1(N890), .IN2(n270), .IN3(N1003), .IN4(n131), .Q(n404) );
  AO221X1 U588 ( .IN1(N439), .IN2(n14), .IN3(N371), .IN4(n348), .IN5(n405), 
        .Q(n402) );
  AO22X1 U589 ( .IN1(N551), .IN2(n124), .IN3(N777), .IN4(n126), .Q(n405) );
  OR4X1 U590 ( .IN1(n406), .IN2(n407), .IN3(n408), .IN4(n409), .Q(N2805) );
  AO221X1 U591 ( .IN1(N2266), .IN2(n329), .IN3(N2611), .IN4(n330), .IN5(n410), 
        .Q(n409) );
  AO22X1 U592 ( .IN1(N292), .IN2(n12), .IN3(N2726), .IN4(n332), .Q(n410) );
  AO222X1 U593 ( .IN1(N2151), .IN2(n333), .IN3(n21), .IN4(n334), .IN5(N1116), 
        .IN6(n335), .Q(n408) );
  AND2X1 U594 ( .IN1(N2381), .IN2(n336), .Q(n407) );
  OA21X1 U595 ( .IN1(n411), .IN2(n412), .IN3(n339), .Q(n406) );
  AO221X1 U596 ( .IN1(N1231), .IN2(n137), .IN3(N1921), .IN4(n340), .IN5(n413), 
        .Q(n412) );
  AO22X1 U597 ( .IN1(N1346), .IN2(n304), .IN3(n21), .IN4(n309), .Q(n413) );
  AO221X1 U598 ( .IN1(N1461), .IN2(n134), .IN3(n342), .IN4(n414), .IN5(n415), 
        .Q(n411) );
  AO22X1 U599 ( .IN1(N1691), .IN2(n85), .IN3(N1806), .IN4(n170), .Q(n415) );
  OR2X1 U600 ( .IN1(n416), .IN2(n417), .Q(n414) );
  AO221X1 U601 ( .IN1(n21), .IN2(n235), .IN3(N1116), .IN4(n129), .IN5(n418), 
        .Q(n417) );
  AO22X1 U602 ( .IN1(N889), .IN2(n270), .IN3(N1002), .IN4(n131), .Q(n418) );
  AO221X1 U603 ( .IN1(N438), .IN2(n14), .IN3(N370), .IN4(n348), .IN5(n419), 
        .Q(n416) );
  AO22X1 U604 ( .IN1(N550), .IN2(n124), .IN3(N776), .IN4(n126), .Q(n419) );
  OR4X1 U605 ( .IN1(n420), .IN2(n421), .IN3(n422), .IN4(n423), .Q(N2804) );
  AO221X1 U606 ( .IN1(n22), .IN2(n329), .IN3(N2610), .IN4(n330), .IN5(n424), 
        .Q(n423) );
  AO22X1 U607 ( .IN1(N291), .IN2(n12), .IN3(n22), .IN4(n332), .Q(n424) );
  AO222X1 U608 ( .IN1(N2150), .IN2(n333), .IN3(n4), .IN4(n334), .IN5(N662), 
        .IN6(n335), .Q(n422) );
  AND2X1 U609 ( .IN1(N2380), .IN2(n336), .Q(n421) );
  OA21X1 U610 ( .IN1(n425), .IN2(n426), .IN3(n339), .Q(n420) );
  AO221X1 U611 ( .IN1(N1230), .IN2(n137), .IN3(N1920), .IN4(n340), .IN5(n427), 
        .Q(n426) );
  AO22X1 U612 ( .IN1(n22), .IN2(n304), .IN3(n4), .IN4(n309), .Q(n427) );
  AO221X1 U613 ( .IN1(N1460), .IN2(n134), .IN3(n342), .IN4(n428), .IN5(n429), 
        .Q(n425) );
  AO22X1 U614 ( .IN1(N1690), .IN2(n85), .IN3(n22), .IN4(n170), .Q(n429) );
  OR2X1 U615 ( .IN1(n430), .IN2(n431), .Q(n428) );
  AO221X1 U616 ( .IN1(n4), .IN2(n235), .IN3(N662), .IN4(n129), .IN5(n432), .Q(
        n431) );
  AO22X1 U617 ( .IN1(n22), .IN2(n270), .IN3(N1001), .IN4(n131), .Q(n432) );
  AO221X1 U618 ( .IN1(n22), .IN2(n14), .IN3(N369), .IN4(n348), .IN5(n433), .Q(
        n430) );
  AO22X1 U619 ( .IN1(N549), .IN2(n124), .IN3(N775), .IN4(n126), .Q(n433) );
  OR4X1 U620 ( .IN1(n434), .IN2(n435), .IN3(n436), .IN4(n437), .Q(N2803) );
  AO221X1 U621 ( .IN1(N436), .IN2(n329), .IN3(n23), .IN4(n330), .IN5(n438), 
        .Q(n437) );
  AO22X1 U622 ( .IN1(N290), .IN2(n12), .IN3(N436), .IN4(n332), .Q(n438) );
  AND2X1 U623 ( .IN1(n63), .IN2(n323), .Q(n332) );
  NAND4X0 U624 ( .IN1(n27), .IN2(n28), .IN3(n29), .IN4(n439), .QN(n323) );
  AO21X1 U625 ( .IN1(n19), .IN2(n440), .IN3(n26), .Q(n439) );
  NOR2X0 U626 ( .IN1(n441), .IN2(n65), .QN(n63) );
  NOR2X0 U627 ( .IN1(n142), .IN2(n65), .QN(n330) );
  AND2X1 U628 ( .IN1(n442), .IN2(n98), .Q(n329) );
  INVX0 U629 ( .INP(n140), .ZN(n98) );
  AO222X1 U630 ( .IN1(n23), .IN2(n333), .IN3(N436), .IN4(n334), .IN5(N436), 
        .IN6(n335), .Q(n436) );
  AND2X1 U631 ( .IN1(n443), .IN2(n89), .Q(n335) );
  INVX0 U632 ( .INP(n83), .ZN(n89) );
  AND2X1 U633 ( .IN1(n442), .IN2(n444), .Q(n334) );
  AND2X1 U634 ( .IN1(n445), .IN2(n90), .Q(n333) );
  INVX0 U635 ( .INP(n152), .ZN(n90) );
  AND2X1 U636 ( .IN1(n23), .IN2(n336), .Q(n435) );
  AND2X1 U637 ( .IN1(n442), .IN2(n99), .Q(n336) );
  OA21X1 U638 ( .IN1(n446), .IN2(n447), .IN3(n339), .Q(n434) );
  AO221X1 U639 ( .IN1(n23), .IN2(n137), .IN3(n23), .IN4(n340), .IN5(n448), .Q(
        n447) );
  AO22X1 U640 ( .IN1(N436), .IN2(n304), .IN3(N436), .IN4(n309), .Q(n448) );
  INVX0 U641 ( .INP(n158), .ZN(n340) );
  AO221X1 U642 ( .IN1(n23), .IN2(n134), .IN3(n342), .IN4(n449), .IN5(n450), 
        .Q(n446) );
  AO22X1 U643 ( .IN1(n23), .IN2(n85), .IN3(N436), .IN4(n170), .Q(n450) );
  INVX0 U644 ( .INP(n73), .ZN(n170) );
  OR2X1 U645 ( .IN1(n451), .IN2(n452), .Q(n449) );
  AO221X1 U646 ( .IN1(N436), .IN2(n235), .IN3(N436), .IN4(n129), .IN5(n453), 
        .Q(n452) );
  AO22X1 U647 ( .IN1(N436), .IN2(n270), .IN3(n23), .IN4(n131), .Q(n453) );
  AO221X1 U648 ( .IN1(N436), .IN2(n14), .IN3(N368), .IN4(n348), .IN5(n454), 
        .Q(n451) );
  AO22X1 U649 ( .IN1(n23), .IN2(n124), .IN3(n23), .IN4(n126), .Q(n454) );
  AND2X1 U650 ( .IN1(n455), .IN2(n145), .Q(n348) );
  NAND3X0 U651 ( .IN1(n106), .IN2(n456), .IN3(n339), .QN(N2802) );
  AND2X1 U652 ( .IN1(n445), .IN2(n152), .Q(n443) );
  AND3X1 U653 ( .IN1(n105), .IN2(n140), .IN3(n442), .Q(n445) );
  AND3X1 U654 ( .IN1(n441), .IN2(n142), .IN3(n13), .Q(n442) );
  MUX21X1 U655 ( .IN1(N264), .IN2(N236), .S(n15), .Q(n65) );
  NAND3X0 U656 ( .IN1(n458), .IN2(n459), .IN3(n460), .QN(n142) );
  NAND2X0 U657 ( .IN1(n461), .IN2(n462), .QN(n458) );
  NAND2X0 U658 ( .IN1(n463), .IN2(n464), .QN(n456) );
  NAND3X0 U659 ( .IN1(n23), .IN2(n465), .IN3(n466), .QN(n464) );
  AND3X1 U660 ( .IN1(n455), .IN2(n175), .IN3(n342), .Q(n106) );
  INVX0 U661 ( .INP(n467), .ZN(n342) );
  NOR4X0 U662 ( .IN1(n468), .IN2(n469), .IN3(n460), .IN4(n322), .QN(N2768) );
  INVX0 U663 ( .INP(n470), .ZN(n460) );
  OR3X1 U664 ( .IN1(n471), .IN2(N2767), .IN3(n472), .Q(n468) );
  NAND4X0 U665 ( .IN1(n473), .IN2(n474), .IN3(n475), .IN4(n476), .QN(N2767) );
  NOR2X0 U666 ( .IN1(n477), .IN2(n478), .QN(n475) );
  NOR4X0 U667 ( .IN1(n479), .IN2(n480), .IN3(n472), .IN4(n481), .QN(N2766) );
  NAND3X0 U668 ( .IN1(n476), .IN2(n482), .IN3(n483), .QN(n479) );
  NOR4X0 U669 ( .IN1(n484), .IN2(n480), .IN3(n485), .IN4(n486), .QN(N2765) );
  NAND4X0 U670 ( .IN1(n441), .IN2(n470), .IN3(n487), .IN4(n474), .QN(n480) );
  AND2X1 U671 ( .IN1(n488), .IN2(n489), .Q(n487) );
  INVX0 U672 ( .INP(n322), .ZN(n441) );
  NOR3X0 U673 ( .IN1(n324), .IN2(n490), .IN3(n141), .QN(n322) );
  NAND3X0 U674 ( .IN1(n105), .IN2(n491), .IN3(n265), .QN(n141) );
  NOR2X0 U675 ( .IN1(n80), .IN2(n281), .QN(n265) );
  NAND3X0 U676 ( .IN1(n310), .IN2(n492), .IN3(n75), .QN(n281) );
  NOR2X0 U677 ( .IN1(n99), .IN2(n444), .QN(n105) );
  INVX0 U678 ( .INP(n123), .ZN(n444) );
  NAND3X0 U679 ( .IN1(n493), .IN2(n459), .IN3(n472), .QN(n123) );
  INVX0 U680 ( .INP(n494), .ZN(n472) );
  NAND2X0 U681 ( .IN1(n461), .IN2(n495), .QN(n493) );
  INVX0 U682 ( .INP(n173), .ZN(n99) );
  NAND3X0 U683 ( .IN1(n496), .IN2(n459), .IN3(n497), .QN(n173) );
  NAND2X0 U684 ( .IN1(n461), .IN2(n21), .QN(n496) );
  NAND3X0 U685 ( .IN1(n470), .IN2(n494), .IN3(n498), .QN(n324) );
  NAND4X0 U686 ( .IN1(n499), .IN2(n500), .IN3(n501), .IN4(n502), .QN(n484) );
  NAND4X0 U687 ( .IN1(n473), .IN2(n470), .IN3(n503), .IN4(n504), .QN(N2764) );
  AND4X1 U688 ( .IN1(n505), .IN2(n506), .IN3(n502), .IN4(n507), .Q(n504) );
  NOR2X0 U689 ( .IN1(n508), .IN2(n497), .QN(n503) );
  INVX0 U690 ( .INP(n483), .ZN(n497) );
  NAND4X0 U691 ( .IN1(n509), .IN2(n498), .IN3(n510), .IN4(n494), .QN(n470) );
  NAND3X0 U692 ( .IN1(n128), .IN2(n510), .IN3(n498), .QN(n494) );
  INVX0 U693 ( .INP(n103), .ZN(n128) );
  NAND2X0 U694 ( .IN1(n491), .IN2(n240), .QN(n103) );
  NOR2X0 U695 ( .IN1(n467), .IN2(n247), .QN(n240) );
  AND4X1 U696 ( .IN1(n474), .IN2(n489), .IN3(n507), .IN4(n511), .Q(n498) );
  NOR2X0 U697 ( .IN1(n512), .IN2(n469), .QN(n511) );
  NAND4X0 U698 ( .IN1(n483), .IN2(n513), .IN3(n499), .IN4(n514), .QN(n469) );
  NAND4X0 U699 ( .IN1(n515), .IN2(n516), .IN3(n517), .IN4(n513), .QN(n483) );
  NOR2X0 U700 ( .IN1(n518), .IN2(n508), .QN(n517) );
  INVX0 U701 ( .INP(n100), .ZN(n515) );
  NAND4X0 U702 ( .IN1(n171), .IN2(n82), .IN3(n152), .IN4(n83), .QN(n100) );
  INVX0 U703 ( .INP(n215), .ZN(n171) );
  NAND3X0 U704 ( .IN1(n519), .IN2(n156), .IN3(n303), .QN(n215) );
  INVX0 U705 ( .INP(n264), .ZN(n303) );
  NAND3X0 U706 ( .IN1(n520), .IN2(n185), .IN3(n521), .QN(n264) );
  INVX0 U707 ( .INP(n122), .ZN(n509) );
  NAND2X0 U708 ( .IN1(n248), .IN2(n491), .QN(n122) );
  INVX0 U709 ( .INP(n95), .ZN(n491) );
  NAND3X0 U710 ( .IN1(n152), .IN2(n83), .IN3(n140), .QN(n95) );
  NAND3X0 U711 ( .IN1(n522), .IN2(n459), .IN3(n485), .QN(n140) );
  INVX0 U712 ( .INP(n513), .ZN(n485) );
  NAND3X0 U713 ( .IN1(n523), .IN2(n152), .IN3(n192), .QN(n513) );
  NOR2X0 U714 ( .IN1(n203), .IN2(n467), .QN(n192) );
  NAND2X0 U715 ( .IN1(n524), .IN2(n492), .QN(n467) );
  NAND3X0 U716 ( .IN1(n525), .IN2(n179), .IN3(n526), .QN(n203) );
  NAND3X0 U717 ( .IN1(n21), .IN2(n527), .IN3(n461), .QN(n522) );
  INVX0 U718 ( .INP(n514), .ZN(n518) );
  NAND3X0 U719 ( .IN1(n23), .IN2(n466), .IN3(n461), .QN(n528) );
  INVX0 U720 ( .INP(n499), .ZN(n508) );
  NAND2X0 U721 ( .IN1(n136), .IN2(n523), .QN(n499) );
  AND2X1 U722 ( .IN1(n516), .IN2(n514), .Q(n523) );
  NAND2X0 U723 ( .IN1(n81), .IN2(n516), .QN(n514) );
  INVX0 U724 ( .INP(n157), .ZN(n81) );
  NAND2X0 U725 ( .IN1(n274), .IN2(n519), .QN(n157) );
  INVX0 U726 ( .INP(n70), .ZN(n519) );
  NAND2X0 U727 ( .IN1(n530), .IN2(n151), .QN(n70) );
  NOR3X0 U728 ( .IN1(n137), .IN2(n283), .IN3(n295), .QN(n274) );
  INVX0 U729 ( .INP(n91), .ZN(n136) );
  NAND2X0 U730 ( .IN1(n524), .IN2(n255), .QN(n91) );
  NOR2X0 U731 ( .IN1(n271), .IN2(n532), .QN(n255) );
  NAND2X0 U732 ( .IN1(n526), .IN2(n533), .QN(n271) );
  INVX0 U733 ( .INP(n534), .ZN(n524) );
  NAND2X0 U734 ( .IN1(n461), .IN2(n466), .QN(n529) );
  NOR4X0 U735 ( .IN1(n9), .IN2(N2037), .IN3(n11), .IN4(a[30]), .QN(n461) );
  NOR2X0 U736 ( .IN1(n262), .IN2(n534), .QN(n248) );
  NAND2X0 U737 ( .IN1(n82), .IN2(n75), .QN(n534) );
  NOR2X0 U738 ( .IN1(n85), .IN2(n309), .QN(n75) );
  INVX0 U739 ( .INP(n151), .ZN(n309) );
  INVX0 U740 ( .INP(n156), .ZN(n85) );
  AO21X1 U741 ( .IN1(n535), .IN2(n536), .IN3(n489), .Q(n156) );
  OR2X1 U742 ( .IN1(n462), .IN2(n19), .Q(n536) );
  INVX0 U743 ( .INP(n80), .ZN(n82) );
  NAND2X0 U744 ( .IN1(n158), .IN2(n73), .QN(n80) );
  AO21X1 U745 ( .IN1(n535), .IN2(n537), .IN3(n474), .Q(n73) );
  OR2X1 U746 ( .IN1(n440), .IN2(n19), .Q(n537) );
  NAND2X0 U747 ( .IN1(n471), .IN2(n459), .QN(n158) );
  INVX0 U748 ( .INP(n507), .ZN(n471) );
  NAND3X0 U749 ( .IN1(n531), .IN2(n474), .IN3(n538), .QN(n507) );
  INVX0 U750 ( .INP(n79), .ZN(n538) );
  NAND3X0 U751 ( .IN1(n266), .IN2(n151), .IN3(n492), .QN(n79) );
  INVX0 U752 ( .INP(n476), .ZN(n541) );
  NAND2X0 U753 ( .IN1(n535), .IN2(n495), .QN(n539) );
  NOR2X0 U754 ( .IN1(n284), .IN2(n129), .QN(n266) );
  MUX21X1 U755 ( .IN1(n542), .IN2(n296), .S(n166), .Q(n284) );
  MUX21X1 U756 ( .IN1(n543), .IN2(n544), .S(n154), .Q(n296) );
  NAND2X0 U757 ( .IN1(n74), .IN2(n531), .QN(n474) );
  INVX0 U758 ( .INP(n155), .ZN(n74) );
  NAND2X0 U759 ( .IN1(n208), .IN2(n205), .QN(n155) );
  NOR3X0 U760 ( .IN1(n304), .IN2(n137), .IN3(n227), .QN(n208) );
  MUX21X1 U761 ( .IN1(n545), .IN2(n272), .S(n182), .Q(n227) );
  MUX21X1 U762 ( .IN1(n543), .IN2(n285), .S(n166), .Q(n272) );
  MUX21X1 U763 ( .IN1(n546), .IN2(n547), .S(n154), .Q(n285) );
  AND3X1 U764 ( .IN1(n510), .IN2(n489), .IN3(n548), .Q(n531) );
  NAND2X0 U765 ( .IN1(n492), .IN2(n308), .QN(n262) );
  INVX0 U766 ( .INP(n532), .ZN(n492) );
  NAND2X0 U767 ( .IN1(n530), .IN2(n185), .QN(n532) );
  NOR2X0 U768 ( .IN1(n134), .IN2(n304), .QN(n530) );
  INVX0 U769 ( .INP(n205), .ZN(n134) );
  AND4X1 U770 ( .IN1(n489), .IN2(n482), .IN3(n501), .IN4(n549), .Q(n473) );
  INVX0 U771 ( .INP(n550), .ZN(n501) );
  NAND3X0 U772 ( .IN1(n172), .IN2(n510), .IN3(n548), .QN(n489) );
  INVX0 U773 ( .INP(n512), .ZN(n548) );
  NAND4X0 U774 ( .IN1(n476), .IN2(n482), .IN3(n551), .IN4(n552), .QN(n512) );
  NOR3X0 U775 ( .IN1(n478), .IN2(n477), .IN3(n550), .QN(n552) );
  INVX0 U776 ( .INP(n500), .ZN(n478) );
  NAND4X0 U777 ( .IN1(n135), .IN2(n553), .IN3(n205), .IN4(n500), .QN(n476) );
  INVX0 U778 ( .INP(n482), .ZN(n555) );
  NAND3X0 U779 ( .IN1(n316), .IN2(n500), .IN3(n553), .QN(n482) );
  INVX0 U780 ( .INP(n556), .ZN(n316) );
  MUX21X1 U781 ( .IN1(n146), .IN2(n557), .S(n304), .Q(n556) );
  INVX0 U782 ( .INP(n147), .ZN(n304) );
  MUX21X1 U783 ( .IN1(n247), .IN2(n184), .S(n185), .Q(n146) );
  MUX21X1 U784 ( .IN1(n558), .IN2(n210), .S(n182), .Q(n184) );
  MUX21X1 U785 ( .IN1(n559), .IN2(n232), .S(n166), .Q(n210) );
  OA222X1 U786 ( .IN1(n560), .IN2(n249), .IN3(n179), .IN4(n561), .IN5(n154), 
        .IN6(n562), .Q(n232) );
  AOI222X1 U787 ( .IN1(n235), .IN2(n563), .IN3(n124), .IN4(n564), .IN5(n236), 
        .IN6(n565), .QN(n249) );
  NAND2X0 U788 ( .IN1(n455), .IN2(n566), .QN(n247) );
  AND2X1 U789 ( .IN1(n521), .IN2(n178), .Q(n455) );
  AND3X1 U790 ( .IN1(n179), .IN2(n149), .IN3(n526), .Q(n521) );
  NOR2X0 U791 ( .IN1(n295), .IN2(n270), .QN(n526) );
  NAND2X0 U792 ( .IN1(n182), .IN2(n166), .QN(n295) );
  NAND2X0 U793 ( .IN1(n535), .IN2(n21), .QN(n554) );
  INVX0 U794 ( .INP(n319), .ZN(n135) );
  MUX21X1 U795 ( .IN1(n302), .IN2(n183), .S(n147), .Q(n319) );
  AO21X1 U796 ( .IN1(n535), .IN2(n567), .IN3(n500), .Q(n147) );
  NAND2X0 U797 ( .IN1(n553), .IN2(n313), .QN(n500) );
  MUX21X1 U798 ( .IN1(n138), .IN2(n520), .S(n137), .Q(n313) );
  INVX0 U799 ( .INP(n568), .ZN(n138) );
  MUX21X1 U800 ( .IN1(n559), .IN2(n181), .S(n182), .Q(n568) );
  MUX21X1 U801 ( .IN1(n209), .IN2(n562), .S(n131), .Q(n181) );
  OA222X1 U802 ( .IN1(n560), .IN2(n229), .IN3(n179), .IN4(n569), .IN5(n154), 
        .IN6(n570), .Q(n209) );
  INVX0 U803 ( .INP(n253), .ZN(n229) );
  AO222X1 U804 ( .IN1(n235), .IN2(n564), .IN3(n124), .IN4(n571), .IN5(n236), 
        .IN6(n572), .Q(n253) );
  NOR2X0 U805 ( .IN1(n573), .IN2(n550), .QN(n553) );
  AO21X1 U806 ( .IN1(n21), .IN2(n527), .IN3(n19), .Q(n567) );
  MUX21X1 U807 ( .IN1(n207), .IN2(n557), .S(n137), .Q(n183) );
  INVX0 U808 ( .INP(n308), .ZN(n557) );
  NOR2X0 U809 ( .IN1(n574), .IN2(n129), .QN(n308) );
  MUX21X1 U810 ( .IN1(n239), .IN2(n546), .S(n129), .Q(n207) );
  MUX21X1 U811 ( .IN1(n250), .IN2(n558), .S(n131), .Q(n239) );
  AOI222X1 U812 ( .IN1(n270), .IN2(n525), .IN3(n126), .IN4(n575), .IN5(n267), 
        .IN6(n269), .QN(n250) );
  INVX0 U813 ( .INP(n69), .ZN(n172) );
  AO21X1 U814 ( .IN1(n137), .IN2(n302), .IN3(n576), .Q(n69) );
  MUX21X1 U815 ( .IN1(n577), .IN2(n574), .S(n129), .Q(n576) );
  OR3X1 U816 ( .IN1(n560), .IN2(n131), .IN3(n543), .Q(n574) );
  AND2X1 U817 ( .IN1(n185), .IN2(n238), .Q(n577) );
  MUX21X1 U818 ( .IN1(n273), .IN2(n546), .S(n131), .Q(n238) );
  OA222X1 U819 ( .IN1(n179), .IN2(n559), .IN3(n154), .IN4(n558), .IN5(n560), 
        .IN6(n578), .Q(n273) );
  INVX0 U820 ( .INP(n525), .ZN(n559) );
  MUX21X1 U821 ( .IN1(n579), .IN2(n580), .S(n149), .Q(n525) );
  INVX0 U822 ( .INP(n310), .ZN(n302) );
  NOR2X0 U823 ( .IN1(n545), .IN2(n129), .QN(n310) );
  INVX0 U824 ( .INP(n182), .ZN(n129) );
  NAND3X0 U825 ( .IN1(n267), .IN2(n166), .IN3(n581), .QN(n545) );
  INVX0 U826 ( .INP(n185), .ZN(n137) );
  NOR2X0 U827 ( .IN1(n573), .IN2(n305), .QN(n550) );
  MUX21X1 U828 ( .IN1(n562), .IN2(n139), .S(n182), .Q(n305) );
  INVX0 U829 ( .INP(n584), .ZN(n477) );
  NAND3X0 U830 ( .IN1(n23), .IN2(n535), .IN3(n466), .QN(n583) );
  MUX21X1 U831 ( .IN1(n283), .IN2(n167), .S(n166), .Q(n139) );
  INVX0 U832 ( .INP(n131), .ZN(n166) );
  NOR2X0 U833 ( .IN1(n549), .IN2(n465), .QN(n131) );
  MUX21X1 U834 ( .IN1(n544), .IN2(n212), .S(n154), .Q(n167) );
  MUX21X1 U835 ( .IN1(n585), .IN2(n231), .S(n179), .Q(n212) );
  AOI222X1 U836 ( .IN1(n235), .IN2(n571), .IN3(n124), .IN4(n586), .IN5(n236), 
        .IN6(n587), .QN(n231) );
  MUX21X1 U837 ( .IN1(n569), .IN2(n546), .S(n126), .Q(n544) );
  INVX0 U838 ( .INP(n566), .ZN(n546) );
  AOI222X1 U839 ( .IN1(n236), .IN2(n563), .IN3(n124), .IN4(n588), .IN5(n235), 
        .IN6(n520), .QN(n569) );
  MUX21X1 U840 ( .IN1(n570), .IN2(n542), .S(n270), .Q(n283) );
  MUX21X1 U841 ( .IN1(n561), .IN2(n543), .S(n126), .Q(n570) );
  NAND2X0 U842 ( .IN1(n589), .IN2(n590), .QN(n543) );
  AOI222X1 U843 ( .IN1(n235), .IN2(n566), .IN3(n124), .IN4(n591), .IN5(n236), 
        .IN6(n592), .QN(n561) );
  INVX0 U844 ( .INP(n533), .ZN(n562) );
  MUX21X1 U845 ( .IN1(n575), .IN2(n581), .S(n126), .Q(n533) );
  INVX0 U846 ( .INP(n542), .ZN(n581) );
  NAND2X0 U847 ( .IN1(n589), .IN2(n579), .QN(n542) );
  NOR2X0 U848 ( .IN1(n593), .IN2(n177), .QN(n589) );
  AO222X1 U849 ( .IN1(n124), .IN2(n566), .IN3(n235), .IN4(n590), .IN5(n236), 
        .IN6(n594), .Q(n575) );
  AO222X1 U850 ( .IN1(n175), .IN2(n193), .IN3(\sub_114_I2_aco/B[0] ), .IN4(
        n320), .IN5(n579), .IN6(n14), .Q(n566) );
  NAND3X0 U851 ( .IN1(n510), .IN2(n584), .IN3(n551), .QN(n573) );
  NAND3X0 U852 ( .IN1(n510), .IN2(n132), .IN3(n551), .QN(n584) );
  AND4X1 U853 ( .IN1(n549), .IN2(n488), .IN3(n595), .IN4(n596), .Q(n551) );
  NOR2X0 U854 ( .IN1(n486), .IN2(n481), .QN(n596) );
  INVX0 U855 ( .INP(n463), .ZN(n595) );
  NOR2X0 U856 ( .IN1(n490), .IN2(n597), .QN(n463) );
  NAND4X0 U857 ( .IN1(n598), .IN2(n599), .IN3(n287), .IN4(n488), .QN(n549) );
  AO222X1 U858 ( .IN1(n270), .IN2(n600), .IN3(n126), .IN4(n269), .IN5(n267), 
        .IN6(n186), .Q(n287) );
  AO222X1 U859 ( .IN1(n235), .IN2(n565), .IN3(n124), .IN4(n572), .IN5(n236), 
        .IN6(n230), .Q(n186) );
  AO222X1 U860 ( .IN1(\sub_114_I2_aco/B[0] ), .IN2(n297), .IN3(n14), .IN4(n306), .IN5(n175), .IN6(n288), .Q(n230) );
  AO222X1 U861 ( .IN1(n235), .IN2(n592), .IN3(n124), .IN4(n563), .IN5(n236), 
        .IN6(n586), .Q(n269) );
  AO222X1 U862 ( .IN1(\sub_114_I2_aco/B[0] ), .IN2(n87), .IN3(n14), .IN4(n92), 
        .IN5(n175), .IN6(n86), .Q(n563) );
  INVX0 U863 ( .INP(n294), .ZN(n132) );
  OA222X1 U864 ( .IN1(n560), .IN2(n168), .IN3(n179), .IN4(n578), .IN5(n154), 
        .IN6(n547), .Q(n294) );
  MUX21X1 U865 ( .IN1(n558), .IN2(n585), .S(n179), .Q(n547) );
  AOI222X1 U866 ( .IN1(n236), .IN2(n564), .IN3(n124), .IN4(n594), .IN5(n235), 
        .IN6(n580), .QN(n585) );
  MUX21X1 U867 ( .IN1(n590), .IN2(n588), .S(n178), .Q(n580) );
  AO222X1 U868 ( .IN1(\sub_114_I2_aco/B[0] ), .IN2(n101), .IN3(n14), .IN4(n193), .IN5(n175), .IN6(n96), .Q(n588) );
  AO222X1 U869 ( .IN1(\sub_114_I2_aco/B[0] ), .IN2(n86), .IN3(n177), .IN4(n87), 
        .IN5(n175), .IN6(n77), .Q(n564) );
  INVX0 U870 ( .INP(n520), .ZN(n558) );
  MUX21X1 U871 ( .IN1(n579), .IN2(n591), .S(n178), .Q(n520) );
  AO222X1 U872 ( .IN1(n175), .IN2(n101), .IN3(\sub_114_I2_aco/B[0] ), .IN4(
        n193), .IN5(n14), .IN6(n590), .Q(n591) );
  MUX21X1 U873 ( .IN1(n601), .IN2(n320), .S(n121), .Q(n590) );
  MUX21X1 U874 ( .IN1(N242), .IN2(N214), .S(n15), .Q(n320) );
  MUX21X1 U875 ( .IN1(N243), .IN2(N215), .S(n15), .Q(n193) );
  AND2X1 U876 ( .IN1(n601), .IN2(n121), .Q(n579) );
  MUX21X1 U877 ( .IN1(N241), .IN2(N213), .S(n15), .Q(n601) );
  INVX0 U878 ( .INP(n600), .ZN(n578) );
  AO222X1 U879 ( .IN1(n235), .IN2(n594), .IN3(n124), .IN4(n592), .IN5(n236), 
        .IN6(n571), .Q(n600) );
  AO222X1 U880 ( .IN1(\sub_114_I2_aco/B[0] ), .IN2(n77), .IN3(n177), .IN4(n86), 
        .IN5(n175), .IN6(n71), .Q(n571) );
  MUX21X1 U881 ( .IN1(N248), .IN2(N220), .S(n15), .Q(n86) );
  AO222X1 U882 ( .IN1(\sub_114_I2_aco/B[0] ), .IN2(n92), .IN3(n177), .IN4(n96), 
        .IN5(n175), .IN6(n87), .Q(n592) );
  MUX21X1 U883 ( .IN1(N247), .IN2(N219), .S(n15), .Q(n87) );
  AO222X1 U884 ( .IN1(\sub_114_I2_aco/B[0] ), .IN2(n96), .IN3(n177), .IN4(n101), .IN5(n175), .IN6(n92), .Q(n594) );
  MUX21X1 U885 ( .IN1(N246), .IN2(N218), .S(n15), .Q(n92) );
  MUX21X1 U886 ( .IN1(N244), .IN2(N216), .S(n15), .Q(n101) );
  MUX21X1 U887 ( .IN1(N245), .IN2(N217), .S(n15), .Q(n96) );
  AOI222X1 U888 ( .IN1(n235), .IN2(n586), .IN3(n124), .IN4(n565), .IN5(n236), 
        .IN6(n234), .QN(n168) );
  AO222X1 U889 ( .IN1(\sub_114_I2_aco/B[0] ), .IN2(n66), .IN3(n177), .IN4(n71), 
        .IN5(n175), .IN6(n317), .Q(n565) );
  AO222X1 U890 ( .IN1(\sub_114_I2_aco/B[0] ), .IN2(n71), .IN3(n177), .IN4(n77), 
        .IN5(n175), .IN6(n66), .Q(n586) );
  MUX21X1 U891 ( .IN1(N249), .IN2(N221), .S(n15), .Q(n77) );
  MUX21X1 U892 ( .IN1(N250), .IN2(N222), .S(n15), .Q(n71) );
  INVX0 U893 ( .INP(n267), .ZN(n560) );
  NOR2X0 U894 ( .IN1(n270), .IN2(n126), .QN(n267) );
  INVX0 U895 ( .INP(n179), .ZN(n126) );
  AO21X1 U896 ( .IN1(n465), .IN2(n462), .IN3(n502), .Q(n179) );
  NAND2X0 U897 ( .IN1(N662), .IN2(N1116), .QN(n462) );
  INVX0 U898 ( .INP(n154), .ZN(n270) );
  AO21X1 U899 ( .IN1(n465), .IN2(n440), .IN3(n488), .Q(n154) );
  NAND3X0 U900 ( .IN1(n599), .IN2(n127), .IN3(n598), .QN(n488) );
  INVX0 U901 ( .INP(n481), .ZN(n598) );
  NAND3X0 U902 ( .IN1(n602), .IN2(n506), .IN3(n502), .QN(n481) );
  NAND4X0 U903 ( .IN1(n599), .IN2(n254), .IN3(n602), .IN4(n506), .QN(n502) );
  AO222X1 U904 ( .IN1(n235), .IN2(n587), .IN3(n124), .IN4(n234), .IN5(n236), 
        .IN6(n187), .Q(n254) );
  AO222X1 U905 ( .IN1(\sub_114_I2_aco/B[0] ), .IN2(n275), .IN3(n177), .IN4(
        n288), .IN5(n175), .IN6(n256), .Q(n187) );
  AO222X1 U906 ( .IN1(\sub_114_I2_aco/B[0] ), .IN2(n306), .IN3(n177), .IN4(
        n314), .IN5(n175), .IN6(n297), .Q(n234) );
  AO222X1 U907 ( .IN1(n235), .IN2(n572), .IN3(n124), .IN4(n587), .IN5(n236), 
        .IN6(n219), .Q(n127) );
  AO222X1 U908 ( .IN1(\sub_114_I2_aco/B[0] ), .IN2(n288), .IN3(n177), .IN4(
        n297), .IN5(n175), .IN6(n275), .Q(n219) );
  MUX21X1 U909 ( .IN1(N255), .IN2(N227), .S(n15), .Q(n297) );
  MUX21X1 U910 ( .IN1(N256), .IN2(N228), .S(n457), .Q(n288) );
  INVX0 U911 ( .INP(n593), .ZN(n236) );
  NAND2X0 U912 ( .IN1(n149), .IN2(n178), .QN(n593) );
  AO222X1 U913 ( .IN1(\sub_114_I2_aco/B[0] ), .IN2(n314), .IN3(n177), .IN4(
        n317), .IN5(n175), .IN6(n306), .Q(n587) );
  MUX21X1 U914 ( .IN1(N254), .IN2(N226), .S(n457), .Q(n306) );
  INVX0 U915 ( .INP(n178), .ZN(n124) );
  AO21X1 U916 ( .IN1(n465), .IN2(n21), .IN3(n506), .Q(n178) );
  AO222X1 U917 ( .IN1(\sub_114_I2_aco/B[0] ), .IN2(n317), .IN3(n177), .IN4(n66), .IN5(n175), .IN6(n314), .Q(n572) );
  MUX21X1 U918 ( .IN1(N253), .IN2(N225), .S(n457), .Q(n314) );
  MUX21X1 U919 ( .IN1(N251), .IN2(N223), .S(n457), .Q(n66) );
  MUX21X1 U920 ( .IN1(N252), .IN2(N224), .S(n457), .Q(n317) );
  INVX0 U921 ( .INP(n149), .ZN(n235) );
  AO21X1 U922 ( .IN1(n465), .IN2(n495), .IN3(n602), .Q(n149) );
  NAND3X0 U923 ( .IN1(n125), .IN2(n506), .IN3(n599), .QN(n602) );
  NAND2X0 U924 ( .IN1(n599), .IN2(n218), .QN(n506) );
  AO222X1 U925 ( .IN1(\sub_114_I2_aco/B[0] ), .IN2(n176), .IN3(n14), .IN4(n256), .IN5(n175), .IN6(n150), .Q(n218) );
  MUX21X1 U926 ( .IN1(N260), .IN2(N232), .S(n457), .Q(n150) );
  AO222X1 U927 ( .IN1(\sub_114_I2_aco/B[0] ), .IN2(n256), .IN3(n14), .IN4(n275), .IN5(n175), .IN6(n176), .Q(n125) );
  MUX21X1 U928 ( .IN1(N259), .IN2(N231), .S(n457), .Q(n176) );
  MUX21X1 U929 ( .IN1(N257), .IN2(N229), .S(n457), .Q(n275) );
  INVX0 U930 ( .INP(n145), .ZN(n177) );
  NAND2X0 U931 ( .IN1(n603), .IN2(n604), .QN(n145) );
  NAND3X0 U932 ( .IN1(n21), .IN2(n527), .IN3(n465), .QN(n604) );
  INVX0 U933 ( .INP(n605), .ZN(n527) );
  INVX0 U934 ( .INP(n606), .ZN(n603) );
  MUX21X1 U935 ( .IN1(N258), .IN2(N230), .S(n457), .Q(n256) );
  AO21X1 U936 ( .IN1(n466), .IN2(n465), .IN3(n505), .Q(n121) );
  AO21X1 U937 ( .IN1(n23), .IN2(n22), .IN3(n21), .Q(n495) );
  NOR3X0 U938 ( .IN1(n109), .IN2(n490), .IN3(n486), .QN(n599) );
  NAND2X0 U939 ( .IN1(n606), .IN2(n505), .QN(n486) );
  NAND4X0 U940 ( .IN1(n597), .IN2(n510), .IN3(n119), .IN4(n505), .QN(n606) );
  NAND3X0 U941 ( .IN1(n597), .IN2(n120), .IN3(n510), .QN(n505) );
  MUX21X1 U942 ( .IN1(N262), .IN2(N234), .S(n457), .Q(n120) );
  MUX21X1 U943 ( .IN1(N261), .IN2(N233), .S(n457), .Q(n119) );
  INVX0 U944 ( .INP(n109), .ZN(n597) );
  INVX0 U945 ( .INP(n510), .ZN(n490) );
  MUX21X1 U946 ( .IN1(N263), .IN2(N235), .S(n457), .Q(n109) );
  AOI22X1 U947 ( .IN1(N59), .IN2(n607), .IN3(N237), .IN4(n608), .QN(n457) );
  NAND2X0 U948 ( .IN1(n605), .IN2(N1116), .QN(n440) );
  NOR2X0 U949 ( .IN1(n23), .IN2(n22), .QN(n605) );
  MUX21X1 U950 ( .IN1(a_in[23]), .IN2(b_in[23]), .S(N54), .Q(N436) );
  INVX0 U951 ( .INP(n540), .ZN(n465) );
  OR2X1 U952 ( .IN1(x[4]), .IN2(x[3]), .Q(n609) );
  NAND2X0 U953 ( .IN1(n535), .IN2(n19), .QN(n540) );
  MUX21X1 U954 ( .IN1(a_in[26]), .IN2(b_in[26]), .S(n36), .Q(N2037) );
  NAND2X0 U955 ( .IN1(n466), .IN2(n535), .QN(n582) );
  INVX0 U956 ( .INP(n459), .ZN(n535) );
  NAND4X0 U957 ( .IN1(n26), .IN2(n27), .IN3(n28), .IN4(n29), .QN(n459) );
  MUX21X1 U958 ( .IN1(a_in[30]), .IN2(b_in[30]), .S(N54), .Q(a[30]) );
  MUX21X1 U959 ( .IN1(a_in[29]), .IN2(b_in[29]), .S(n36), .Q(a[29]) );
  MUX21X1 U960 ( .IN1(a_in[28]), .IN2(b_in[28]), .S(n36), .Q(a[28]) );
  MUX21X1 U961 ( .IN1(a_in[27]), .IN2(b_in[27]), .S(N54), .Q(a[27]) );
  NOR2X0 U962 ( .IN1(N1116), .IN2(N662), .QN(n466) );
  MUX21X1 U963 ( .IN1(a_in[24]), .IN2(b_in[24]), .S(n36), .Q(N662) );
  MUX21X1 U964 ( .IN1(a_in[25]), .IN2(b_in[25]), .S(n36), .Q(N1116) );
  AO222X1 U965 ( .IN1(N140), .IN2(n18), .IN3(N164), .IN4(n608), .IN5(N188), 
        .IN6(n607), .Q(N236) );
  AO222X1 U966 ( .IN1(N139), .IN2(n18), .IN3(N163), .IN4(n608), .IN5(N187), 
        .IN6(n607), .Q(N235) );
  AO222X1 U967 ( .IN1(N138), .IN2(n18), .IN3(N162), .IN4(n608), .IN5(N186), 
        .IN6(n607), .Q(N234) );
  AO222X1 U968 ( .IN1(N137), .IN2(n18), .IN3(N161), .IN4(n608), .IN5(N185), 
        .IN6(n607), .Q(N233) );
  AO222X1 U969 ( .IN1(N136), .IN2(n18), .IN3(N160), .IN4(n608), .IN5(N184), 
        .IN6(n607), .Q(N232) );
  AO222X1 U970 ( .IN1(N135), .IN2(n18), .IN3(N159), .IN4(n608), .IN5(N183), 
        .IN6(n607), .Q(N231) );
  AO222X1 U971 ( .IN1(N134), .IN2(n18), .IN3(N158), .IN4(n608), .IN5(N182), 
        .IN6(n607), .Q(N230) );
  AO222X1 U972 ( .IN1(N133), .IN2(n18), .IN3(N157), .IN4(n608), .IN5(N181), 
        .IN6(n607), .Q(N229) );
  AO222X1 U973 ( .IN1(N132), .IN2(n18), .IN3(N156), .IN4(n608), .IN5(N180), 
        .IN6(n607), .Q(N228) );
  AO222X1 U974 ( .IN1(N131), .IN2(n18), .IN3(N155), .IN4(n608), .IN5(N179), 
        .IN6(n607), .Q(N227) );
  AO222X1 U975 ( .IN1(N130), .IN2(n18), .IN3(N154), .IN4(n17), .IN5(N178), 
        .IN6(n16), .Q(N226) );
  AO222X1 U976 ( .IN1(N129), .IN2(n18), .IN3(N153), .IN4(n608), .IN5(N177), 
        .IN6(n607), .Q(N225) );
  AO222X1 U977 ( .IN1(N128), .IN2(n610), .IN3(N152), .IN4(n17), .IN5(N176), 
        .IN6(n16), .Q(N224) );
  AO222X1 U978 ( .IN1(N127), .IN2(n610), .IN3(N151), .IN4(n17), .IN5(N175), 
        .IN6(n16), .Q(N223) );
  AO222X1 U979 ( .IN1(N126), .IN2(n610), .IN3(N150), .IN4(n17), .IN5(N174), 
        .IN6(n16), .Q(N222) );
  AO222X1 U980 ( .IN1(N125), .IN2(n610), .IN3(N149), .IN4(n17), .IN5(N173), 
        .IN6(n16), .Q(N221) );
  AO222X1 U981 ( .IN1(N124), .IN2(n610), .IN3(N148), .IN4(n17), .IN5(N172), 
        .IN6(n16), .Q(N220) );
  AO222X1 U982 ( .IN1(N123), .IN2(n610), .IN3(N147), .IN4(n17), .IN5(N171), 
        .IN6(n16), .Q(N219) );
  AO222X1 U983 ( .IN1(N122), .IN2(n610), .IN3(N146), .IN4(n17), .IN5(N170), 
        .IN6(n16), .Q(N218) );
  AO222X1 U984 ( .IN1(N121), .IN2(n610), .IN3(N145), .IN4(n17), .IN5(N169), 
        .IN6(n16), .Q(N217) );
  AO222X1 U985 ( .IN1(N120), .IN2(n610), .IN3(N144), .IN4(n17), .IN5(N168), 
        .IN6(n16), .Q(N216) );
  AO222X1 U986 ( .IN1(N119), .IN2(n610), .IN3(N143), .IN4(n17), .IN5(N167), 
        .IN6(n16), .Q(N215) );
  AO222X1 U987 ( .IN1(N118), .IN2(n610), .IN3(N142), .IN4(n17), .IN5(N166), 
        .IN6(n16), .Q(N214) );
  AO222X1 U988 ( .IN1(N117), .IN2(n18), .IN3(N141), .IN4(n17), .IN5(N165), 
        .IN6(n16), .Q(N213) );
  XNOR2X1 U989 ( .IN1(n25), .IN2(n31), .Q(n610) );
  MUX21X1 U990 ( .IN1(a_in[31]), .IN2(b_in[31]), .S(n36), .Q(a[31]) );
  MUX21X1 U991 ( .IN1(b_in[31]), .IN2(a_in[31]), .S(n36), .Q(b[31]) );
endmodule


module fpalu_multiplier_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[8]), .IN2(A[8]), .Q(SUM[8]) );
endmodule


module fpalu_multiplier_DW01_inc_1 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(SUM[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module fpalu_multiplier_DW01_add_1 ( A, B, CI, SUM, CO );
  input [45:0] A;
  input [45:0] B;
  output [45:0] SUM;
  input CI;
  output CO;
  wire   \A[22] , \A[21] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104;
  assign SUM[22] = \A[22] ;
  assign \A[22]  = A[22];
  assign SUM[21] = \A[21] ;
  assign \A[21]  = A[21];

  INVX0 U2 ( .INP(n26), .ZN(n2) );
  INVX0 U3 ( .INP(n98), .ZN(n20) );
  INVX0 U4 ( .INP(n93), .ZN(n19) );
  INVX0 U5 ( .INP(n89), .ZN(n18) );
  INVX0 U6 ( .INP(n86), .ZN(n17) );
  INVX0 U7 ( .INP(n82), .ZN(n16) );
  INVX0 U8 ( .INP(n78), .ZN(n15) );
  INVX0 U9 ( .INP(n74), .ZN(n14) );
  INVX0 U10 ( .INP(n70), .ZN(n13) );
  INVX0 U11 ( .INP(n66), .ZN(n12) );
  INVX0 U12 ( .INP(n62), .ZN(n11) );
  INVX0 U13 ( .INP(n58), .ZN(n10) );
  INVX0 U14 ( .INP(n54), .ZN(n9) );
  INVX0 U15 ( .INP(n50), .ZN(n8) );
  INVX0 U16 ( .INP(n46), .ZN(n7) );
  INVX0 U17 ( .INP(n42), .ZN(n6) );
  INVX0 U18 ( .INP(n38), .ZN(n5) );
  INVX0 U19 ( .INP(n34), .ZN(n4) );
  INVX0 U20 ( .INP(n30), .ZN(n3) );
  INVX0 U21 ( .INP(n102), .ZN(n21) );
  AND2X1 U22 ( .IN1(n101), .IN2(n1), .Q(SUM[23]) );
  OR2X1 U23 ( .IN1(B[23]), .IN2(A[23]), .Q(n1) );
  XNOR2X1 U24 ( .IN1(n22), .IN2(B[45]), .Q(SUM[45]) );
  AOI22X1 U25 ( .IN1(n23), .IN2(B[44]), .IN3(n24), .IN4(A[44]), .QN(n22) );
  OR2X1 U26 ( .IN1(A[44]), .IN2(n24), .Q(n23) );
  XOR3X1 U27 ( .IN1(B[44]), .IN2(A[44]), .IN3(n24), .Q(SUM[44]) );
  OAI21X1 U28 ( .IN1(n25), .IN2(n26), .IN3(n27), .QN(n24) );
  XOR2X1 U29 ( .IN1(n28), .IN2(n25), .Q(SUM[43]) );
  OA21X1 U30 ( .IN1(n29), .IN2(n30), .IN3(n31), .Q(n25) );
  NAND2X0 U31 ( .IN1(n2), .IN2(n27), .QN(n28) );
  NAND2X0 U32 ( .IN1(B[43]), .IN2(A[43]), .QN(n27) );
  NOR2X0 U33 ( .IN1(B[43]), .IN2(A[43]), .QN(n26) );
  XOR2X1 U34 ( .IN1(n32), .IN2(n29), .Q(SUM[42]) );
  OA21X1 U35 ( .IN1(n33), .IN2(n34), .IN3(n35), .Q(n29) );
  NAND2X0 U36 ( .IN1(n3), .IN2(n31), .QN(n32) );
  NAND2X0 U37 ( .IN1(B[42]), .IN2(A[42]), .QN(n31) );
  NOR2X0 U38 ( .IN1(B[42]), .IN2(A[42]), .QN(n30) );
  XOR2X1 U39 ( .IN1(n36), .IN2(n33), .Q(SUM[41]) );
  OA21X1 U40 ( .IN1(n37), .IN2(n38), .IN3(n39), .Q(n33) );
  NAND2X0 U41 ( .IN1(n4), .IN2(n35), .QN(n36) );
  NAND2X0 U42 ( .IN1(B[41]), .IN2(A[41]), .QN(n35) );
  NOR2X0 U43 ( .IN1(B[41]), .IN2(A[41]), .QN(n34) );
  XOR2X1 U44 ( .IN1(n40), .IN2(n37), .Q(SUM[40]) );
  OA21X1 U45 ( .IN1(n41), .IN2(n42), .IN3(n43), .Q(n37) );
  NAND2X0 U46 ( .IN1(n5), .IN2(n39), .QN(n40) );
  NAND2X0 U47 ( .IN1(B[40]), .IN2(A[40]), .QN(n39) );
  NOR2X0 U48 ( .IN1(B[40]), .IN2(A[40]), .QN(n38) );
  XOR2X1 U49 ( .IN1(n44), .IN2(n41), .Q(SUM[39]) );
  OA21X1 U50 ( .IN1(n45), .IN2(n46), .IN3(n47), .Q(n41) );
  NAND2X0 U51 ( .IN1(n6), .IN2(n43), .QN(n44) );
  NAND2X0 U52 ( .IN1(B[39]), .IN2(A[39]), .QN(n43) );
  NOR2X0 U53 ( .IN1(B[39]), .IN2(A[39]), .QN(n42) );
  XOR2X1 U54 ( .IN1(n48), .IN2(n45), .Q(SUM[38]) );
  OA21X1 U55 ( .IN1(n49), .IN2(n50), .IN3(n51), .Q(n45) );
  NAND2X0 U56 ( .IN1(n7), .IN2(n47), .QN(n48) );
  NAND2X0 U57 ( .IN1(B[38]), .IN2(A[38]), .QN(n47) );
  NOR2X0 U58 ( .IN1(B[38]), .IN2(A[38]), .QN(n46) );
  XOR2X1 U59 ( .IN1(n52), .IN2(n49), .Q(SUM[37]) );
  OA21X1 U60 ( .IN1(n53), .IN2(n54), .IN3(n55), .Q(n49) );
  NAND2X0 U61 ( .IN1(n8), .IN2(n51), .QN(n52) );
  NAND2X0 U62 ( .IN1(B[37]), .IN2(A[37]), .QN(n51) );
  NOR2X0 U63 ( .IN1(B[37]), .IN2(A[37]), .QN(n50) );
  XOR2X1 U64 ( .IN1(n56), .IN2(n53), .Q(SUM[36]) );
  OA21X1 U65 ( .IN1(n57), .IN2(n58), .IN3(n59), .Q(n53) );
  NAND2X0 U66 ( .IN1(n9), .IN2(n55), .QN(n56) );
  NAND2X0 U67 ( .IN1(B[36]), .IN2(A[36]), .QN(n55) );
  NOR2X0 U68 ( .IN1(B[36]), .IN2(A[36]), .QN(n54) );
  XOR2X1 U69 ( .IN1(n60), .IN2(n57), .Q(SUM[35]) );
  OA21X1 U70 ( .IN1(n61), .IN2(n62), .IN3(n63), .Q(n57) );
  NAND2X0 U71 ( .IN1(n10), .IN2(n59), .QN(n60) );
  NAND2X0 U72 ( .IN1(B[35]), .IN2(A[35]), .QN(n59) );
  NOR2X0 U73 ( .IN1(B[35]), .IN2(A[35]), .QN(n58) );
  XOR2X1 U74 ( .IN1(n64), .IN2(n61), .Q(SUM[34]) );
  OA21X1 U75 ( .IN1(n65), .IN2(n66), .IN3(n67), .Q(n61) );
  NAND2X0 U76 ( .IN1(n11), .IN2(n63), .QN(n64) );
  NAND2X0 U77 ( .IN1(B[34]), .IN2(A[34]), .QN(n63) );
  NOR2X0 U78 ( .IN1(B[34]), .IN2(A[34]), .QN(n62) );
  XOR2X1 U79 ( .IN1(n68), .IN2(n65), .Q(SUM[33]) );
  OA21X1 U80 ( .IN1(n69), .IN2(n70), .IN3(n71), .Q(n65) );
  NAND2X0 U81 ( .IN1(n12), .IN2(n67), .QN(n68) );
  NAND2X0 U82 ( .IN1(B[33]), .IN2(A[33]), .QN(n67) );
  NOR2X0 U83 ( .IN1(B[33]), .IN2(A[33]), .QN(n66) );
  XOR2X1 U84 ( .IN1(n72), .IN2(n69), .Q(SUM[32]) );
  OA21X1 U85 ( .IN1(n73), .IN2(n74), .IN3(n75), .Q(n69) );
  NAND2X0 U86 ( .IN1(n13), .IN2(n71), .QN(n72) );
  NAND2X0 U87 ( .IN1(B[32]), .IN2(A[32]), .QN(n71) );
  NOR2X0 U88 ( .IN1(B[32]), .IN2(A[32]), .QN(n70) );
  XOR2X1 U89 ( .IN1(n76), .IN2(n73), .Q(SUM[31]) );
  OA21X1 U90 ( .IN1(n77), .IN2(n78), .IN3(n79), .Q(n73) );
  NAND2X0 U91 ( .IN1(n14), .IN2(n75), .QN(n76) );
  NAND2X0 U92 ( .IN1(B[31]), .IN2(A[31]), .QN(n75) );
  NOR2X0 U93 ( .IN1(B[31]), .IN2(A[31]), .QN(n74) );
  XOR2X1 U94 ( .IN1(n80), .IN2(n77), .Q(SUM[30]) );
  OA21X1 U95 ( .IN1(n81), .IN2(n82), .IN3(n83), .Q(n77) );
  NAND2X0 U96 ( .IN1(n15), .IN2(n79), .QN(n80) );
  NAND2X0 U97 ( .IN1(B[30]), .IN2(A[30]), .QN(n79) );
  NOR2X0 U98 ( .IN1(B[30]), .IN2(A[30]), .QN(n78) );
  XOR2X1 U99 ( .IN1(n84), .IN2(n81), .Q(SUM[29]) );
  OA21X1 U100 ( .IN1(n85), .IN2(n86), .IN3(n87), .Q(n81) );
  NAND2X0 U101 ( .IN1(n16), .IN2(n83), .QN(n84) );
  NAND2X0 U102 ( .IN1(B[29]), .IN2(A[29]), .QN(n83) );
  NOR2X0 U103 ( .IN1(B[29]), .IN2(A[29]), .QN(n82) );
  XOR2X1 U104 ( .IN1(n88), .IN2(n85), .Q(SUM[28]) );
  OA21X1 U105 ( .IN1(n89), .IN2(n90), .IN3(n91), .Q(n85) );
  NAND2X0 U106 ( .IN1(n17), .IN2(n87), .QN(n88) );
  NAND2X0 U107 ( .IN1(B[28]), .IN2(A[28]), .QN(n87) );
  NOR2X0 U108 ( .IN1(B[28]), .IN2(A[28]), .QN(n86) );
  XOR2X1 U109 ( .IN1(n92), .IN2(n90), .Q(SUM[27]) );
  OA21X1 U110 ( .IN1(n93), .IN2(n94), .IN3(n95), .Q(n90) );
  NAND2X0 U111 ( .IN1(n18), .IN2(n91), .QN(n92) );
  NAND2X0 U112 ( .IN1(B[27]), .IN2(A[27]), .QN(n91) );
  NOR2X0 U113 ( .IN1(B[27]), .IN2(A[27]), .QN(n89) );
  XOR2X1 U114 ( .IN1(n96), .IN2(n94), .Q(SUM[26]) );
  OA21X1 U115 ( .IN1(n97), .IN2(n98), .IN3(n99), .Q(n94) );
  NAND2X0 U116 ( .IN1(n19), .IN2(n95), .QN(n96) );
  NAND2X0 U117 ( .IN1(B[26]), .IN2(A[26]), .QN(n95) );
  NOR2X0 U118 ( .IN1(B[26]), .IN2(A[26]), .QN(n93) );
  XOR2X1 U119 ( .IN1(n100), .IN2(n97), .Q(SUM[25]) );
  OA21X1 U120 ( .IN1(n101), .IN2(n102), .IN3(n103), .Q(n97) );
  NAND2X0 U121 ( .IN1(n20), .IN2(n99), .QN(n100) );
  NAND2X0 U122 ( .IN1(B[25]), .IN2(A[25]), .QN(n99) );
  NOR2X0 U123 ( .IN1(B[25]), .IN2(A[25]), .QN(n98) );
  XOR2X1 U124 ( .IN1(n104), .IN2(n101), .Q(SUM[24]) );
  NAND2X0 U125 ( .IN1(n21), .IN2(n103), .QN(n104) );
  NAND2X0 U126 ( .IN1(B[24]), .IN2(A[24]), .QN(n103) );
  NOR2X0 U127 ( .IN1(B[24]), .IN2(A[24]), .QN(n102) );
  NAND2X0 U128 ( .IN1(B[23]), .IN2(A[23]), .QN(n101) );
endmodule


module fpalu_multiplier_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [23:0] A;
  input [23:0] B;
  output [47:0] PRODUCT;
  input TC;
  wire   \ab[23][23] , \ab[23][22] , \ab[23][21] , \ab[23][20] , \ab[23][19] ,
         \ab[23][18] , \ab[23][17] , \ab[23][16] , \ab[23][15] , \ab[23][14] ,
         \ab[23][13] , \ab[23][12] , \ab[23][11] , \ab[23][10] , \ab[23][9] ,
         \ab[23][8] , \ab[23][7] , \ab[23][6] , \ab[23][5] , \ab[23][4] ,
         \ab[23][3] , \ab[23][2] , \ab[23][1] , \ab[23][0] , \ab[22][23] ,
         \ab[22][22] , \ab[22][21] , \ab[22][20] , \ab[22][19] , \ab[22][18] ,
         \ab[22][17] , \ab[22][16] , \ab[22][15] , \ab[22][14] , \ab[22][13] ,
         \ab[22][12] , \ab[22][11] , \ab[22][10] , \ab[22][9] , \ab[22][8] ,
         \ab[22][7] , \ab[22][6] , \ab[22][5] , \ab[22][4] , \ab[22][3] ,
         \ab[22][2] , \ab[22][1] , \ab[22][0] , \ab[21][23] , \ab[21][22] ,
         \ab[21][21] , \ab[21][20] , \ab[21][19] , \ab[21][18] , \ab[21][17] ,
         \ab[21][16] , \ab[21][15] , \ab[21][14] , \ab[21][13] , \ab[21][12] ,
         \ab[21][11] , \ab[21][10] , \ab[21][9] , \ab[21][8] , \ab[21][7] ,
         \ab[21][6] , \ab[21][5] , \ab[21][4] , \ab[21][3] , \ab[21][2] ,
         \ab[21][1] , \ab[21][0] , \ab[20][23] , \ab[20][22] , \ab[20][21] ,
         \ab[20][20] , \ab[20][19] , \ab[20][18] , \ab[20][17] , \ab[20][16] ,
         \ab[20][15] , \ab[20][14] , \ab[20][13] , \ab[20][12] , \ab[20][11] ,
         \ab[20][10] , \ab[20][9] , \ab[20][8] , \ab[20][7] , \ab[20][6] ,
         \ab[20][5] , \ab[20][4] , \ab[20][3] , \ab[20][2] , \ab[20][1] ,
         \ab[20][0] , \ab[19][23] , \ab[19][22] , \ab[19][21] , \ab[19][20] ,
         \ab[19][19] , \ab[19][18] , \ab[19][17] , \ab[19][16] , \ab[19][15] ,
         \ab[19][14] , \ab[19][13] , \ab[19][12] , \ab[19][11] , \ab[19][10] ,
         \ab[19][9] , \ab[19][8] , \ab[19][7] , \ab[19][6] , \ab[19][5] ,
         \ab[19][4] , \ab[19][3] , \ab[19][2] , \ab[19][1] , \ab[19][0] ,
         \ab[18][23] , \ab[18][22] , \ab[18][21] , \ab[18][20] , \ab[18][19] ,
         \ab[18][18] , \ab[18][17] , \ab[18][16] , \ab[18][15] , \ab[18][14] ,
         \ab[18][13] , \ab[18][12] , \ab[18][11] , \ab[18][10] , \ab[18][9] ,
         \ab[18][8] , \ab[18][7] , \ab[18][6] , \ab[18][5] , \ab[18][4] ,
         \ab[18][3] , \ab[18][2] , \ab[18][1] , \ab[18][0] , \ab[17][23] ,
         \ab[17][22] , \ab[17][21] , \ab[17][20] , \ab[17][19] , \ab[17][18] ,
         \ab[17][17] , \ab[17][16] , \ab[17][15] , \ab[17][14] , \ab[17][13] ,
         \ab[17][12] , \ab[17][11] , \ab[17][10] , \ab[17][9] , \ab[17][8] ,
         \ab[17][7] , \ab[17][6] , \ab[17][5] , \ab[17][4] , \ab[17][3] ,
         \ab[17][2] , \ab[17][1] , \ab[17][0] , \ab[16][23] , \ab[16][22] ,
         \ab[16][21] , \ab[16][20] , \ab[16][19] , \ab[16][18] , \ab[16][17] ,
         \ab[16][16] , \ab[16][15] , \ab[16][14] , \ab[16][13] , \ab[16][12] ,
         \ab[16][11] , \ab[16][10] , \ab[16][9] , \ab[16][8] , \ab[16][7] ,
         \ab[16][6] , \ab[16][5] , \ab[16][4] , \ab[16][3] , \ab[16][2] ,
         \ab[16][1] , \ab[16][0] , \ab[15][23] , \ab[15][22] , \ab[15][21] ,
         \ab[15][20] , \ab[15][19] , \ab[15][18] , \ab[15][17] , \ab[15][16] ,
         \ab[15][15] , \ab[15][14] , \ab[15][13] , \ab[15][12] , \ab[15][11] ,
         \ab[15][10] , \ab[15][9] , \ab[15][8] , \ab[15][7] , \ab[15][6] ,
         \ab[15][5] , \ab[15][4] , \ab[15][3] , \ab[15][2] , \ab[15][1] ,
         \ab[15][0] , \ab[14][23] , \ab[14][22] , \ab[14][21] , \ab[14][20] ,
         \ab[14][19] , \ab[14][18] , \ab[14][17] , \ab[14][16] , \ab[14][15] ,
         \ab[14][14] , \ab[14][13] , \ab[14][12] , \ab[14][11] , \ab[14][10] ,
         \ab[14][9] , \ab[14][8] , \ab[14][7] , \ab[14][6] , \ab[14][5] ,
         \ab[14][4] , \ab[14][3] , \ab[14][2] , \ab[14][1] , \ab[14][0] ,
         \ab[13][23] , \ab[13][22] , \ab[13][21] , \ab[13][20] , \ab[13][19] ,
         \ab[13][18] , \ab[13][17] , \ab[13][16] , \ab[13][15] , \ab[13][14] ,
         \ab[13][13] , \ab[13][12] , \ab[13][11] , \ab[13][10] , \ab[13][9] ,
         \ab[13][8] , \ab[13][7] , \ab[13][6] , \ab[13][5] , \ab[13][4] ,
         \ab[13][3] , \ab[13][2] , \ab[13][1] , \ab[13][0] , \ab[12][23] ,
         \ab[12][22] , \ab[12][21] , \ab[12][20] , \ab[12][19] , \ab[12][18] ,
         \ab[12][17] , \ab[12][16] , \ab[12][15] , \ab[12][14] , \ab[12][13] ,
         \ab[12][12] , \ab[12][11] , \ab[12][10] , \ab[12][9] , \ab[12][8] ,
         \ab[12][7] , \ab[12][6] , \ab[12][5] , \ab[12][4] , \ab[12][3] ,
         \ab[12][2] , \ab[12][1] , \ab[12][0] , \ab[11][23] , \ab[11][22] ,
         \ab[11][21] , \ab[11][20] , \ab[11][19] , \ab[11][18] , \ab[11][17] ,
         \ab[11][16] , \ab[11][15] , \ab[11][14] , \ab[11][13] , \ab[11][12] ,
         \ab[11][11] , \ab[11][10] , \ab[11][9] , \ab[11][8] , \ab[11][7] ,
         \ab[11][6] , \ab[11][5] , \ab[11][4] , \ab[11][3] , \ab[11][2] ,
         \ab[11][1] , \ab[11][0] , \ab[10][23] , \ab[10][22] , \ab[10][21] ,
         \ab[10][20] , \ab[10][19] , \ab[10][18] , \ab[10][17] , \ab[10][16] ,
         \ab[10][15] , \ab[10][14] , \ab[10][13] , \ab[10][12] , \ab[10][11] ,
         \ab[10][10] , \ab[10][9] , \ab[10][8] , \ab[10][7] , \ab[10][6] ,
         \ab[10][5] , \ab[10][4] , \ab[10][3] , \ab[10][2] , \ab[10][1] ,
         \ab[10][0] , \ab[9][23] , \ab[9][22] , \ab[9][21] , \ab[9][20] ,
         \ab[9][19] , \ab[9][18] , \ab[9][17] , \ab[9][16] , \ab[9][15] ,
         \ab[9][14] , \ab[9][13] , \ab[9][12] , \ab[9][11] , \ab[9][10] ,
         \ab[9][9] , \ab[9][8] , \ab[9][7] , \ab[9][6] , \ab[9][5] ,
         \ab[9][4] , \ab[9][3] , \ab[9][2] , \ab[9][1] , \ab[9][0] ,
         \ab[8][23] , \ab[8][22] , \ab[8][21] , \ab[8][20] , \ab[8][19] ,
         \ab[8][18] , \ab[8][17] , \ab[8][16] , \ab[8][15] , \ab[8][14] ,
         \ab[8][13] , \ab[8][12] , \ab[8][11] , \ab[8][10] , \ab[8][9] ,
         \ab[8][8] , \ab[8][7] , \ab[8][6] , \ab[8][5] , \ab[8][4] ,
         \ab[8][3] , \ab[8][2] , \ab[8][1] , \ab[8][0] , \ab[7][23] ,
         \ab[7][22] , \ab[7][21] , \ab[7][20] , \ab[7][19] , \ab[7][18] ,
         \ab[7][17] , \ab[7][16] , \ab[7][15] , \ab[7][14] , \ab[7][13] ,
         \ab[7][12] , \ab[7][11] , \ab[7][10] , \ab[7][9] , \ab[7][8] ,
         \ab[7][7] , \ab[7][6] , \ab[7][5] , \ab[7][4] , \ab[7][3] ,
         \ab[7][2] , \ab[7][1] , \ab[7][0] , \ab[6][23] , \ab[6][22] ,
         \ab[6][21] , \ab[6][20] , \ab[6][19] , \ab[6][18] , \ab[6][17] ,
         \ab[6][16] , \ab[6][15] , \ab[6][14] , \ab[6][13] , \ab[6][12] ,
         \ab[6][11] , \ab[6][10] , \ab[6][9] , \ab[6][8] , \ab[6][7] ,
         \ab[6][6] , \ab[6][5] , \ab[6][4] , \ab[6][3] , \ab[6][2] ,
         \ab[6][1] , \ab[6][0] , \ab[5][23] , \ab[5][22] , \ab[5][21] ,
         \ab[5][20] , \ab[5][19] , \ab[5][18] , \ab[5][17] , \ab[5][16] ,
         \ab[5][15] , \ab[5][14] , \ab[5][13] , \ab[5][12] , \ab[5][11] ,
         \ab[5][10] , \ab[5][9] , \ab[5][8] , \ab[5][7] , \ab[5][6] ,
         \ab[5][5] , \ab[5][4] , \ab[5][3] , \ab[5][2] , \ab[5][1] ,
         \ab[5][0] , \ab[4][23] , \ab[4][22] , \ab[4][21] , \ab[4][20] ,
         \ab[4][19] , \ab[4][18] , \ab[4][17] , \ab[4][16] , \ab[4][15] ,
         \ab[4][14] , \ab[4][13] , \ab[4][12] , \ab[4][11] , \ab[4][10] ,
         \ab[4][9] , \ab[4][8] , \ab[4][7] , \ab[4][6] , \ab[4][5] ,
         \ab[4][4] , \ab[4][3] , \ab[4][2] , \ab[4][1] , \ab[4][0] ,
         \ab[3][23] , \ab[3][22] , \ab[3][21] , \ab[3][20] , \ab[3][19] ,
         \ab[3][18] , \ab[3][17] , \ab[3][16] , \ab[3][15] , \ab[3][14] ,
         \ab[3][13] , \ab[3][12] , \ab[3][11] , \ab[3][10] , \ab[3][9] ,
         \ab[3][8] , \ab[3][7] , \ab[3][6] , \ab[3][5] , \ab[3][4] ,
         \ab[3][3] , \ab[3][2] , \ab[3][1] , \ab[3][0] , \ab[2][23] ,
         \ab[2][22] , \ab[2][21] , \ab[2][20] , \ab[2][19] , \ab[2][18] ,
         \ab[2][17] , \ab[2][16] , \ab[2][15] , \ab[2][14] , \ab[2][13] ,
         \ab[2][12] , \ab[2][11] , \ab[2][10] , \ab[2][9] , \ab[2][8] ,
         \ab[2][7] , \ab[2][6] , \ab[2][5] , \ab[2][4] , \ab[2][3] ,
         \ab[2][2] , \ab[2][1] , \ab[2][0] , \ab[1][23] , \ab[1][22] ,
         \ab[1][21] , \ab[1][20] , \ab[1][19] , \ab[1][18] , \ab[1][17] ,
         \ab[1][16] , \ab[1][15] , \ab[1][14] , \ab[1][13] , \ab[1][12] ,
         \ab[1][11] , \ab[1][10] , \ab[1][9] , \ab[1][8] , \ab[1][7] ,
         \ab[1][6] , \ab[1][5] , \ab[1][4] , \ab[1][3] , \ab[1][2] ,
         \ab[1][1] , \ab[0][23] , \ab[0][22] , \ab[0][21] , \ab[0][20] ,
         \ab[0][19] , \ab[0][18] , \ab[0][17] , \ab[0][16] , \ab[0][15] ,
         \ab[0][14] , \ab[0][13] , \ab[0][12] , \ab[0][11] , \ab[0][10] ,
         \ab[0][9] , \ab[0][8] , \ab[0][7] , \ab[0][6] , \ab[0][5] ,
         \ab[0][4] , \ab[0][3] , \ab[0][2] , \CARRYB[23][22] ,
         \CARRYB[23][21] , \CARRYB[23][20] , \CARRYB[23][19] ,
         \CARRYB[23][18] , \CARRYB[23][17] , \CARRYB[23][16] ,
         \CARRYB[23][15] , \CARRYB[23][14] , \CARRYB[23][13] ,
         \CARRYB[23][12] , \CARRYB[23][11] , \CARRYB[23][10] , \CARRYB[23][9] ,
         \CARRYB[23][8] , \CARRYB[23][7] , \CARRYB[23][6] , \CARRYB[23][5] ,
         \CARRYB[23][4] , \CARRYB[23][3] , \CARRYB[23][2] , \CARRYB[23][1] ,
         \CARRYB[23][0] , \CARRYB[22][22] , \CARRYB[22][21] , \CARRYB[22][20] ,
         \CARRYB[22][19] , \CARRYB[22][18] , \CARRYB[22][17] ,
         \CARRYB[22][16] , \CARRYB[22][15] , \CARRYB[22][14] ,
         \CARRYB[22][13] , \CARRYB[22][12] , \CARRYB[22][11] ,
         \CARRYB[22][10] , \CARRYB[22][9] , \CARRYB[22][8] , \CARRYB[22][7] ,
         \CARRYB[22][6] , \CARRYB[22][5] , \CARRYB[22][4] , \CARRYB[22][3] ,
         \CARRYB[22][2] , \CARRYB[22][1] , \CARRYB[22][0] , \CARRYB[21][22] ,
         \CARRYB[21][21] , \CARRYB[21][20] , \CARRYB[21][19] ,
         \CARRYB[21][18] , \CARRYB[21][17] , \CARRYB[21][16] ,
         \CARRYB[21][15] , \CARRYB[21][14] , \CARRYB[21][13] ,
         \CARRYB[21][12] , \CARRYB[21][11] , \CARRYB[21][10] , \CARRYB[21][9] ,
         \CARRYB[21][8] , \CARRYB[21][7] , \CARRYB[21][6] , \CARRYB[21][5] ,
         \CARRYB[21][4] , \CARRYB[21][3] , \CARRYB[21][2] , \CARRYB[21][1] ,
         \CARRYB[21][0] , \CARRYB[20][22] , \CARRYB[20][21] , \CARRYB[20][20] ,
         \CARRYB[20][19] , \CARRYB[20][18] , \CARRYB[20][17] ,
         \CARRYB[20][16] , \CARRYB[20][15] , \CARRYB[20][14] ,
         \CARRYB[20][13] , \CARRYB[20][12] , \CARRYB[20][11] ,
         \CARRYB[20][10] , \CARRYB[20][9] , \CARRYB[20][8] , \CARRYB[20][7] ,
         \CARRYB[20][6] , \CARRYB[20][5] , \CARRYB[20][4] , \CARRYB[20][3] ,
         \CARRYB[20][2] , \CARRYB[20][1] , \CARRYB[20][0] , \CARRYB[19][22] ,
         \CARRYB[19][21] , \CARRYB[19][20] , \CARRYB[19][19] ,
         \CARRYB[19][18] , \CARRYB[19][17] , \CARRYB[19][16] ,
         \CARRYB[19][15] , \CARRYB[19][14] , \CARRYB[19][13] ,
         \CARRYB[19][12] , \CARRYB[19][11] , \CARRYB[19][10] , \CARRYB[19][9] ,
         \CARRYB[19][8] , \CARRYB[19][7] , \CARRYB[19][6] , \CARRYB[19][5] ,
         \CARRYB[19][4] , \CARRYB[19][3] , \CARRYB[19][2] , \CARRYB[19][1] ,
         \CARRYB[19][0] , \CARRYB[18][22] , \CARRYB[18][21] , \CARRYB[18][20] ,
         \CARRYB[18][19] , \CARRYB[18][18] , \CARRYB[18][17] ,
         \CARRYB[18][16] , \CARRYB[18][15] , \CARRYB[18][14] ,
         \CARRYB[18][13] , \CARRYB[18][12] , \CARRYB[18][11] ,
         \CARRYB[18][10] , \CARRYB[18][9] , \CARRYB[18][8] , \CARRYB[18][7] ,
         \CARRYB[18][6] , \CARRYB[18][5] , \CARRYB[18][4] , \CARRYB[18][3] ,
         \CARRYB[18][2] , \CARRYB[18][1] , \CARRYB[18][0] , \CARRYB[17][22] ,
         \CARRYB[17][21] , \CARRYB[17][20] , \CARRYB[17][19] ,
         \CARRYB[17][18] , \CARRYB[17][17] , \CARRYB[17][16] ,
         \CARRYB[17][15] , \CARRYB[17][14] , \CARRYB[17][13] ,
         \CARRYB[17][12] , \CARRYB[17][11] , \CARRYB[17][10] , \CARRYB[17][9] ,
         \CARRYB[17][8] , \CARRYB[17][7] , \CARRYB[17][6] , \CARRYB[17][5] ,
         \CARRYB[17][4] , \CARRYB[17][3] , \CARRYB[17][2] , \CARRYB[17][1] ,
         \CARRYB[17][0] , \CARRYB[16][22] , \CARRYB[16][21] , \CARRYB[16][20] ,
         \CARRYB[16][19] , \CARRYB[16][18] , \CARRYB[16][17] ,
         \CARRYB[16][16] , \CARRYB[16][15] , \CARRYB[16][14] ,
         \CARRYB[16][13] , \CARRYB[16][12] , \CARRYB[16][11] ,
         \CARRYB[16][10] , \CARRYB[16][9] , \CARRYB[16][8] , \CARRYB[16][7] ,
         \CARRYB[16][6] , \CARRYB[16][5] , \CARRYB[16][4] , \CARRYB[16][3] ,
         \CARRYB[16][2] , \CARRYB[16][1] , \CARRYB[16][0] , \CARRYB[15][22] ,
         \CARRYB[15][21] , \CARRYB[15][20] , \CARRYB[15][19] ,
         \CARRYB[15][18] , \CARRYB[15][17] , \CARRYB[15][16] ,
         \CARRYB[15][15] , \CARRYB[15][14] , \CARRYB[15][13] ,
         \CARRYB[15][12] , \CARRYB[15][11] , \CARRYB[15][10] , \CARRYB[15][9] ,
         \CARRYB[15][8] , \CARRYB[15][7] , \CARRYB[15][6] , \CARRYB[15][5] ,
         \CARRYB[15][4] , \CARRYB[15][3] , \CARRYB[15][2] , \CARRYB[15][1] ,
         \CARRYB[15][0] , \CARRYB[14][22] , \CARRYB[14][21] , \CARRYB[14][20] ,
         \CARRYB[14][19] , \CARRYB[14][18] , \CARRYB[14][17] ,
         \CARRYB[14][16] , \CARRYB[14][15] , \CARRYB[14][14] ,
         \CARRYB[14][13] , \CARRYB[14][12] , \CARRYB[14][11] ,
         \CARRYB[14][10] , \CARRYB[14][9] , \CARRYB[14][8] , \CARRYB[14][7] ,
         \CARRYB[14][6] , \CARRYB[14][5] , \CARRYB[14][4] , \CARRYB[14][3] ,
         \CARRYB[14][2] , \CARRYB[14][1] , \CARRYB[14][0] , \CARRYB[13][22] ,
         \CARRYB[13][21] , \CARRYB[13][20] , \CARRYB[13][19] ,
         \CARRYB[13][18] , \CARRYB[13][17] , \CARRYB[13][16] ,
         \CARRYB[13][15] , \CARRYB[13][14] , \CARRYB[13][13] ,
         \CARRYB[13][12] , \CARRYB[13][11] , \CARRYB[13][10] , \CARRYB[13][9] ,
         \CARRYB[13][8] , \CARRYB[13][7] , \CARRYB[13][6] , \CARRYB[13][5] ,
         \CARRYB[13][4] , \CARRYB[13][3] , \CARRYB[13][2] , \CARRYB[13][1] ,
         \CARRYB[13][0] , \CARRYB[12][22] , \CARRYB[12][21] , \CARRYB[12][20] ,
         \CARRYB[12][19] , \CARRYB[12][18] , \CARRYB[12][17] ,
         \CARRYB[12][16] , \CARRYB[12][15] , \CARRYB[12][14] ,
         \CARRYB[12][13] , \CARRYB[12][12] , \CARRYB[12][11] ,
         \CARRYB[12][10] , \CARRYB[12][9] , \CARRYB[12][8] , \CARRYB[12][7] ,
         \CARRYB[12][6] , \CARRYB[12][5] , \CARRYB[12][4] , \CARRYB[12][3] ,
         \CARRYB[12][2] , \CARRYB[12][1] , \CARRYB[12][0] , \CARRYB[11][22] ,
         \CARRYB[11][21] , \CARRYB[11][20] , \CARRYB[11][19] ,
         \CARRYB[11][18] , \CARRYB[11][17] , \CARRYB[11][16] ,
         \CARRYB[11][15] , \CARRYB[11][14] , \CARRYB[11][13] ,
         \CARRYB[11][12] , \CARRYB[11][11] , \CARRYB[11][10] , \CARRYB[11][9] ,
         \CARRYB[11][8] , \CARRYB[11][7] , \CARRYB[11][6] , \CARRYB[11][5] ,
         \CARRYB[11][4] , \CARRYB[11][3] , \CARRYB[11][2] , \CARRYB[11][1] ,
         \CARRYB[11][0] , \CARRYB[10][22] , \CARRYB[10][21] , \CARRYB[10][20] ,
         \CARRYB[10][19] , \CARRYB[10][18] , \CARRYB[10][17] ,
         \CARRYB[10][16] , \CARRYB[10][15] , \CARRYB[10][14] ,
         \CARRYB[10][13] , \CARRYB[10][12] , \CARRYB[10][11] ,
         \CARRYB[10][10] , \CARRYB[10][9] , \CARRYB[10][8] , \CARRYB[10][7] ,
         \CARRYB[10][6] , \CARRYB[10][5] , \CARRYB[10][4] , \CARRYB[10][3] ,
         \CARRYB[10][2] , \CARRYB[10][1] , \CARRYB[10][0] , \CARRYB[9][22] ,
         \CARRYB[9][21] , \CARRYB[9][20] , \CARRYB[9][19] , \CARRYB[9][18] ,
         \CARRYB[9][17] , \CARRYB[9][16] , \CARRYB[9][15] , \CARRYB[9][14] ,
         \CARRYB[9][13] , \CARRYB[9][12] , \CARRYB[9][11] , \CARRYB[9][10] ,
         \CARRYB[9][9] , \CARRYB[9][8] , \CARRYB[9][7] , \CARRYB[9][6] ,
         \CARRYB[9][5] , \CARRYB[9][4] , \CARRYB[9][3] , \CARRYB[9][2] ,
         \CARRYB[9][1] , \CARRYB[9][0] , \CARRYB[8][22] , \CARRYB[8][21] ,
         \CARRYB[8][20] , \CARRYB[8][19] , \CARRYB[8][18] , \CARRYB[8][17] ,
         \CARRYB[8][16] , \CARRYB[8][15] , \CARRYB[8][14] , \CARRYB[8][13] ,
         \CARRYB[8][12] , \CARRYB[8][11] , \CARRYB[8][10] , \CARRYB[8][9] ,
         \CARRYB[8][8] , \CARRYB[8][7] , \CARRYB[8][6] , \CARRYB[8][5] ,
         \CARRYB[8][4] , \CARRYB[8][3] , \CARRYB[8][2] , \CARRYB[8][1] ,
         \CARRYB[8][0] , \CARRYB[7][22] , \CARRYB[7][21] , \CARRYB[7][20] ,
         \CARRYB[7][19] , \CARRYB[7][18] , \CARRYB[7][17] , \CARRYB[7][16] ,
         \CARRYB[7][15] , \CARRYB[7][14] , \CARRYB[7][13] , \CARRYB[7][12] ,
         \CARRYB[7][11] , \CARRYB[7][10] , \CARRYB[7][9] , \CARRYB[7][8] ,
         \CARRYB[7][7] , \CARRYB[7][6] , \CARRYB[7][5] , \CARRYB[7][4] ,
         \CARRYB[7][3] , \CARRYB[7][2] , \CARRYB[7][1] , \CARRYB[7][0] ,
         \CARRYB[6][22] , \CARRYB[6][21] , \CARRYB[6][20] , \CARRYB[6][19] ,
         \CARRYB[6][18] , \CARRYB[6][17] , \CARRYB[6][16] , \CARRYB[6][15] ,
         \CARRYB[6][14] , \CARRYB[6][13] , \CARRYB[6][12] , \CARRYB[6][11] ,
         \CARRYB[6][10] , \CARRYB[6][9] , \CARRYB[6][8] , \CARRYB[6][7] ,
         \CARRYB[6][6] , \CARRYB[6][5] , \CARRYB[6][4] , \CARRYB[6][3] ,
         \CARRYB[6][2] , \CARRYB[6][1] , \CARRYB[6][0] , \CARRYB[5][22] ,
         \CARRYB[5][21] , \CARRYB[5][20] , \CARRYB[5][19] , \CARRYB[5][18] ,
         \CARRYB[5][17] , \CARRYB[5][16] , \CARRYB[5][15] , \CARRYB[5][14] ,
         \CARRYB[5][13] , \CARRYB[5][12] , \CARRYB[5][11] , \CARRYB[5][10] ,
         \CARRYB[5][9] , \CARRYB[5][8] , \CARRYB[5][7] , \CARRYB[5][6] ,
         \CARRYB[5][5] , \CARRYB[5][4] , \CARRYB[5][3] , \CARRYB[5][2] ,
         \CARRYB[5][1] , \CARRYB[5][0] , \CARRYB[4][22] , \CARRYB[4][21] ,
         \CARRYB[4][20] , \CARRYB[4][19] , \CARRYB[4][18] , \CARRYB[4][17] ,
         \CARRYB[4][16] , \CARRYB[4][15] , \CARRYB[4][14] , \CARRYB[4][13] ,
         \CARRYB[4][12] , \CARRYB[4][11] , \CARRYB[4][10] , \CARRYB[4][9] ,
         \CARRYB[4][8] , \CARRYB[4][7] , \CARRYB[4][6] , \CARRYB[4][5] ,
         \CARRYB[4][4] , \CARRYB[4][3] , \CARRYB[4][2] , \CARRYB[4][1] ,
         \CARRYB[4][0] , \CARRYB[3][22] , \CARRYB[3][21] , \CARRYB[3][20] ,
         \CARRYB[3][19] , \CARRYB[3][18] , \CARRYB[3][17] , \CARRYB[3][16] ,
         \CARRYB[3][15] , \CARRYB[3][14] , \CARRYB[3][13] , \CARRYB[3][12] ,
         \CARRYB[3][11] , \CARRYB[3][10] , \CARRYB[3][9] , \CARRYB[3][8] ,
         \CARRYB[3][7] , \CARRYB[3][6] , \CARRYB[3][5] , \CARRYB[3][4] ,
         \CARRYB[3][3] , \CARRYB[3][2] , \CARRYB[3][1] , \CARRYB[3][0] ,
         \CARRYB[2][22] , \CARRYB[2][21] , \CARRYB[2][20] , \CARRYB[2][19] ,
         \CARRYB[2][18] , \CARRYB[2][17] , \CARRYB[2][16] , \CARRYB[2][15] ,
         \CARRYB[2][14] , \CARRYB[2][13] , \CARRYB[2][12] , \CARRYB[2][11] ,
         \CARRYB[2][10] , \CARRYB[2][9] , \CARRYB[2][8] , \CARRYB[2][7] ,
         \CARRYB[2][6] , \CARRYB[2][5] , \CARRYB[2][4] , \CARRYB[2][3] ,
         \CARRYB[2][2] , \CARRYB[2][1] , \CARRYB[2][0] , \CARRYB[1][0] ,
         \SUMB[23][22] , \SUMB[23][21] , \SUMB[23][20] , \SUMB[23][19] ,
         \SUMB[23][18] , \SUMB[23][17] , \SUMB[23][16] , \SUMB[23][15] ,
         \SUMB[23][14] , \SUMB[23][13] , \SUMB[23][12] , \SUMB[23][11] ,
         \SUMB[23][10] , \SUMB[23][9] , \SUMB[23][8] , \SUMB[23][7] ,
         \SUMB[23][6] , \SUMB[23][5] , \SUMB[23][4] , \SUMB[23][3] ,
         \SUMB[23][2] , \SUMB[23][1] , \SUMB[23][0] , \SUMB[22][22] ,
         \SUMB[22][21] , \SUMB[22][20] , \SUMB[22][19] , \SUMB[22][18] ,
         \SUMB[22][17] , \SUMB[22][16] , \SUMB[22][15] , \SUMB[22][14] ,
         \SUMB[22][13] , \SUMB[22][12] , \SUMB[22][11] , \SUMB[22][10] ,
         \SUMB[22][9] , \SUMB[22][8] , \SUMB[22][7] , \SUMB[22][6] ,
         \SUMB[22][5] , \SUMB[22][4] , \SUMB[22][3] , \SUMB[22][2] ,
         \SUMB[22][1] , \SUMB[21][22] , \SUMB[21][21] , \SUMB[21][20] ,
         \SUMB[21][19] , \SUMB[21][18] , \SUMB[21][17] , \SUMB[21][16] ,
         \SUMB[21][15] , \SUMB[21][14] , \SUMB[21][13] , \SUMB[21][12] ,
         \SUMB[21][11] , \SUMB[21][10] , \SUMB[21][9] , \SUMB[21][8] ,
         \SUMB[21][7] , \SUMB[21][6] , \SUMB[21][5] , \SUMB[21][4] ,
         \SUMB[21][3] , \SUMB[21][2] , \SUMB[21][1] , \SUMB[20][22] ,
         \SUMB[20][21] , \SUMB[20][20] , \SUMB[20][19] , \SUMB[20][18] ,
         \SUMB[20][17] , \SUMB[20][16] , \SUMB[20][15] , \SUMB[20][14] ,
         \SUMB[20][13] , \SUMB[20][12] , \SUMB[20][11] , \SUMB[20][10] ,
         \SUMB[20][9] , \SUMB[20][8] , \SUMB[20][7] , \SUMB[20][6] ,
         \SUMB[20][5] , \SUMB[20][4] , \SUMB[20][3] , \SUMB[20][2] ,
         \SUMB[20][1] , \SUMB[19][22] , \SUMB[19][21] , \SUMB[19][20] ,
         \SUMB[19][19] , \SUMB[19][18] , \SUMB[19][17] , \SUMB[19][16] ,
         \SUMB[19][15] , \SUMB[19][14] , \SUMB[19][13] , \SUMB[19][12] ,
         \SUMB[19][11] , \SUMB[19][10] , \SUMB[19][9] , \SUMB[19][8] ,
         \SUMB[19][7] , \SUMB[19][6] , \SUMB[19][5] , \SUMB[19][4] ,
         \SUMB[19][3] , \SUMB[19][2] , \SUMB[19][1] , \SUMB[18][22] ,
         \SUMB[18][21] , \SUMB[18][20] , \SUMB[18][19] , \SUMB[18][18] ,
         \SUMB[18][17] , \SUMB[18][16] , \SUMB[18][15] , \SUMB[18][14] ,
         \SUMB[18][13] , \SUMB[18][12] , \SUMB[18][11] , \SUMB[18][10] ,
         \SUMB[18][9] , \SUMB[18][8] , \SUMB[18][7] , \SUMB[18][6] ,
         \SUMB[18][5] , \SUMB[18][4] , \SUMB[18][3] , \SUMB[18][2] ,
         \SUMB[18][1] , \SUMB[17][22] , \SUMB[17][21] , \SUMB[17][20] ,
         \SUMB[17][19] , \SUMB[17][18] , \SUMB[17][17] , \SUMB[17][16] ,
         \SUMB[17][15] , \SUMB[17][14] , \SUMB[17][13] , \SUMB[17][12] ,
         \SUMB[17][11] , \SUMB[17][10] , \SUMB[17][9] , \SUMB[17][8] ,
         \SUMB[17][7] , \SUMB[17][6] , \SUMB[17][5] , \SUMB[17][4] ,
         \SUMB[17][3] , \SUMB[17][2] , \SUMB[17][1] , \SUMB[16][22] ,
         \SUMB[16][21] , \SUMB[16][20] , \SUMB[16][19] , \SUMB[16][18] ,
         \SUMB[16][17] , \SUMB[16][16] , \SUMB[16][15] , \SUMB[16][14] ,
         \SUMB[16][13] , \SUMB[16][12] , \SUMB[16][11] , \SUMB[16][10] ,
         \SUMB[16][9] , \SUMB[16][8] , \SUMB[16][7] , \SUMB[16][6] ,
         \SUMB[16][5] , \SUMB[16][4] , \SUMB[16][3] , \SUMB[16][2] ,
         \SUMB[16][1] , \SUMB[15][22] , \SUMB[15][21] , \SUMB[15][20] ,
         \SUMB[15][19] , \SUMB[15][18] , \SUMB[15][17] , \SUMB[15][16] ,
         \SUMB[15][15] , \SUMB[15][14] , \SUMB[15][13] , \SUMB[15][12] ,
         \SUMB[15][11] , \SUMB[15][10] , \SUMB[15][9] , \SUMB[15][8] ,
         \SUMB[15][7] , \SUMB[15][6] , \SUMB[15][5] , \SUMB[15][4] ,
         \SUMB[15][3] , \SUMB[15][2] , \SUMB[15][1] , \SUMB[14][22] ,
         \SUMB[14][21] , \SUMB[14][20] , \SUMB[14][19] , \SUMB[14][18] ,
         \SUMB[14][17] , \SUMB[14][16] , \SUMB[14][15] , \SUMB[14][14] ,
         \SUMB[14][13] , \SUMB[14][12] , \SUMB[14][11] , \SUMB[14][10] ,
         \SUMB[14][9] , \SUMB[14][8] , \SUMB[14][7] , \SUMB[14][6] ,
         \SUMB[14][5] , \SUMB[14][4] , \SUMB[14][3] , \SUMB[14][2] ,
         \SUMB[14][1] , \SUMB[13][22] , \SUMB[13][21] , \SUMB[13][20] ,
         \SUMB[13][19] , \SUMB[13][18] , \SUMB[13][17] , \SUMB[13][16] ,
         \SUMB[13][15] , \SUMB[13][14] , \SUMB[13][13] , \SUMB[13][12] ,
         \SUMB[13][11] , \SUMB[13][10] , \SUMB[13][9] , \SUMB[13][8] ,
         \SUMB[13][7] , \SUMB[13][6] , \SUMB[13][5] , \SUMB[13][4] ,
         \SUMB[13][3] , \SUMB[13][2] , \SUMB[13][1] , \SUMB[12][22] ,
         \SUMB[12][21] , \SUMB[12][20] , \SUMB[12][19] , \SUMB[12][18] ,
         \SUMB[12][17] , \SUMB[12][16] , \SUMB[12][15] , \SUMB[12][14] ,
         \SUMB[12][13] , \SUMB[12][12] , \SUMB[12][11] , \SUMB[12][10] ,
         \SUMB[12][9] , \SUMB[12][8] , \SUMB[12][7] , \SUMB[12][6] ,
         \SUMB[12][5] , \SUMB[12][4] , \SUMB[12][3] , \SUMB[12][2] ,
         \SUMB[12][1] , \SUMB[11][22] , \SUMB[11][21] , \SUMB[11][20] ,
         \SUMB[11][19] , \SUMB[11][18] , \SUMB[11][17] , \SUMB[11][16] ,
         \SUMB[11][15] , \SUMB[11][14] , \SUMB[11][13] , \SUMB[11][12] ,
         \SUMB[11][11] , \SUMB[11][10] , \SUMB[11][9] , \SUMB[11][8] ,
         \SUMB[11][7] , \SUMB[11][6] , \SUMB[11][5] , \SUMB[11][4] ,
         \SUMB[11][3] , \SUMB[11][2] , \SUMB[11][1] , \SUMB[10][22] ,
         \SUMB[10][21] , \SUMB[10][20] , \SUMB[10][19] , \SUMB[10][18] ,
         \SUMB[10][17] , \SUMB[10][16] , \SUMB[10][15] , \SUMB[10][14] ,
         \SUMB[10][13] , \SUMB[10][12] , \SUMB[10][11] , \SUMB[10][10] ,
         \SUMB[10][9] , \SUMB[10][8] , \SUMB[10][7] , \SUMB[10][6] ,
         \SUMB[10][5] , \SUMB[10][4] , \SUMB[10][3] , \SUMB[10][2] ,
         \SUMB[10][1] , \SUMB[9][22] , \SUMB[9][21] , \SUMB[9][20] ,
         \SUMB[9][19] , \SUMB[9][18] , \SUMB[9][17] , \SUMB[9][16] ,
         \SUMB[9][15] , \SUMB[9][14] , \SUMB[9][13] , \SUMB[9][12] ,
         \SUMB[9][11] , \SUMB[9][10] , \SUMB[9][9] , \SUMB[9][8] ,
         \SUMB[9][7] , \SUMB[9][6] , \SUMB[9][5] , \SUMB[9][4] , \SUMB[9][3] ,
         \SUMB[9][2] , \SUMB[9][1] , \SUMB[8][22] , \SUMB[8][21] ,
         \SUMB[8][20] , \SUMB[8][19] , \SUMB[8][18] , \SUMB[8][17] ,
         \SUMB[8][16] , \SUMB[8][15] , \SUMB[8][14] , \SUMB[8][13] ,
         \SUMB[8][12] , \SUMB[8][11] , \SUMB[8][10] , \SUMB[8][9] ,
         \SUMB[8][8] , \SUMB[8][7] , \SUMB[8][6] , \SUMB[8][5] , \SUMB[8][4] ,
         \SUMB[8][3] , \SUMB[8][2] , \SUMB[8][1] , \SUMB[7][22] ,
         \SUMB[7][21] , \SUMB[7][20] , \SUMB[7][19] , \SUMB[7][18] ,
         \SUMB[7][17] , \SUMB[7][16] , \SUMB[7][15] , \SUMB[7][14] ,
         \SUMB[7][13] , \SUMB[7][12] , \SUMB[7][11] , \SUMB[7][10] ,
         \SUMB[7][9] , \SUMB[7][8] , \SUMB[7][7] , \SUMB[7][6] , \SUMB[7][5] ,
         \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] , \SUMB[6][22] ,
         \SUMB[6][21] , \SUMB[6][20] , \SUMB[6][19] , \SUMB[6][18] ,
         \SUMB[6][17] , \SUMB[6][16] , \SUMB[6][15] , \SUMB[6][14] ,
         \SUMB[6][13] , \SUMB[6][12] , \SUMB[6][11] , \SUMB[6][10] ,
         \SUMB[6][9] , \SUMB[6][8] , \SUMB[6][7] , \SUMB[6][6] , \SUMB[6][5] ,
         \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] , \SUMB[5][22] ,
         \SUMB[5][21] , \SUMB[5][20] , \SUMB[5][19] , \SUMB[5][18] ,
         \SUMB[5][17] , \SUMB[5][16] , \SUMB[5][15] , \SUMB[5][14] ,
         \SUMB[5][13] , \SUMB[5][12] , \SUMB[5][11] , \SUMB[5][10] ,
         \SUMB[5][9] , \SUMB[5][8] , \SUMB[5][7] , \SUMB[5][6] , \SUMB[5][5] ,
         \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][22] ,
         \SUMB[4][21] , \SUMB[4][20] , \SUMB[4][19] , \SUMB[4][18] ,
         \SUMB[4][17] , \SUMB[4][16] , \SUMB[4][15] , \SUMB[4][14] ,
         \SUMB[4][13] , \SUMB[4][12] , \SUMB[4][11] , \SUMB[4][10] ,
         \SUMB[4][9] , \SUMB[4][8] , \SUMB[4][7] , \SUMB[4][6] , \SUMB[4][5] ,
         \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][22] ,
         \SUMB[3][21] , \SUMB[3][20] , \SUMB[3][19] , \SUMB[3][18] ,
         \SUMB[3][17] , \SUMB[3][16] , \SUMB[3][15] , \SUMB[3][14] ,
         \SUMB[3][13] , \SUMB[3][12] , \SUMB[3][11] , \SUMB[3][10] ,
         \SUMB[3][9] , \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][22] ,
         \SUMB[2][21] , \SUMB[2][20] , \SUMB[2][19] , \SUMB[2][18] ,
         \SUMB[2][17] , \SUMB[2][16] , \SUMB[2][15] , \SUMB[2][14] ,
         \SUMB[2][13] , \SUMB[2][12] , \SUMB[2][11] , \SUMB[2][10] ,
         \SUMB[2][9] , \SUMB[2][8] , \SUMB[2][7] , \SUMB[2][6] , \SUMB[2][5] ,
         \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] , \SUMB[1][22] ,
         \SUMB[1][21] , \SUMB[1][20] , \SUMB[1][19] , \SUMB[1][18] ,
         \SUMB[1][17] , \SUMB[1][16] , \SUMB[1][15] , \SUMB[1][14] ,
         \SUMB[1][13] , \SUMB[1][12] , \SUMB[1][11] , \SUMB[1][10] ,
         \SUMB[1][9] , \SUMB[1][8] , \SUMB[1][7] , \SUMB[1][6] , \SUMB[1][5] ,
         \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] , \SUMB[1][1] , \A1[44] ,
         \A1[43] , \A1[42] , \A1[41] , \A1[40] , \A1[39] , \A1[38] , \A1[37] ,
         \A1[36] , \A1[35] , \A1[34] , \A1[33] , \A1[32] , \A1[31] , \A1[30] ,
         \A1[29] , \A1[28] , \A1[27] , \A1[26] , \A1[25] , \A1[24] , \A1[23] ,
         \A1[22] , \A1[20] , \A1[19] , \A1[18] , \A1[17] , \A1[16] , \A1[15] ,
         \A1[14] , \A1[13] , \A1[12] , \A1[11] , \A1[10] , \A1[9] , \A1[8] ,
         \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] ,
         \A1[0] , n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
         n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20;
  assign \ab[23][23]  = B[23];

  FADDX1 S4_0 ( .A(\ab[23][0] ), .B(\CARRYB[22][0] ), .CI(\SUMB[22][1] ), .CO(
        \CARRYB[23][0] ), .S(\SUMB[23][0] ) );
  FADDX1 S4_1 ( .A(\ab[23][1] ), .B(\CARRYB[22][1] ), .CI(\SUMB[22][2] ), .CO(
        \CARRYB[23][1] ), .S(\SUMB[23][1] ) );
  FADDX1 S4_2 ( .A(\ab[23][2] ), .B(\CARRYB[22][2] ), .CI(\SUMB[22][3] ), .CO(
        \CARRYB[23][2] ), .S(\SUMB[23][2] ) );
  FADDX1 S4_3 ( .A(\ab[23][3] ), .B(\CARRYB[22][3] ), .CI(\SUMB[22][4] ), .CO(
        \CARRYB[23][3] ), .S(\SUMB[23][3] ) );
  FADDX1 S4_4 ( .A(\ab[23][4] ), .B(\CARRYB[22][4] ), .CI(\SUMB[22][5] ), .CO(
        \CARRYB[23][4] ), .S(\SUMB[23][4] ) );
  FADDX1 S4_5 ( .A(\ab[23][5] ), .B(\CARRYB[22][5] ), .CI(\SUMB[22][6] ), .CO(
        \CARRYB[23][5] ), .S(\SUMB[23][5] ) );
  FADDX1 S4_6 ( .A(\ab[23][6] ), .B(\CARRYB[22][6] ), .CI(\SUMB[22][7] ), .CO(
        \CARRYB[23][6] ), .S(\SUMB[23][6] ) );
  FADDX1 S4_7 ( .A(\ab[23][7] ), .B(\CARRYB[22][7] ), .CI(\SUMB[22][8] ), .CO(
        \CARRYB[23][7] ), .S(\SUMB[23][7] ) );
  FADDX1 S4_8 ( .A(\ab[23][8] ), .B(\CARRYB[22][8] ), .CI(\SUMB[22][9] ), .CO(
        \CARRYB[23][8] ), .S(\SUMB[23][8] ) );
  FADDX1 S4_9 ( .A(\ab[23][9] ), .B(\CARRYB[22][9] ), .CI(\SUMB[22][10] ), 
        .CO(\CARRYB[23][9] ), .S(\SUMB[23][9] ) );
  FADDX1 S4_10 ( .A(\ab[23][10] ), .B(\CARRYB[22][10] ), .CI(\SUMB[22][11] ), 
        .CO(\CARRYB[23][10] ), .S(\SUMB[23][10] ) );
  FADDX1 S4_11 ( .A(\ab[23][11] ), .B(\CARRYB[22][11] ), .CI(\SUMB[22][12] ), 
        .CO(\CARRYB[23][11] ), .S(\SUMB[23][11] ) );
  FADDX1 S4_12 ( .A(\ab[23][12] ), .B(\CARRYB[22][12] ), .CI(\SUMB[22][13] ), 
        .CO(\CARRYB[23][12] ), .S(\SUMB[23][12] ) );
  FADDX1 S4_13 ( .A(\ab[23][13] ), .B(\CARRYB[22][13] ), .CI(\SUMB[22][14] ), 
        .CO(\CARRYB[23][13] ), .S(\SUMB[23][13] ) );
  FADDX1 S4_14 ( .A(\ab[23][14] ), .B(\CARRYB[22][14] ), .CI(\SUMB[22][15] ), 
        .CO(\CARRYB[23][14] ), .S(\SUMB[23][14] ) );
  FADDX1 S4_15 ( .A(\ab[23][15] ), .B(\CARRYB[22][15] ), .CI(\SUMB[22][16] ), 
        .CO(\CARRYB[23][15] ), .S(\SUMB[23][15] ) );
  FADDX1 S4_16 ( .A(\ab[23][16] ), .B(\CARRYB[22][16] ), .CI(\SUMB[22][17] ), 
        .CO(\CARRYB[23][16] ), .S(\SUMB[23][16] ) );
  FADDX1 S4_17 ( .A(\ab[23][17] ), .B(\CARRYB[22][17] ), .CI(\SUMB[22][18] ), 
        .CO(\CARRYB[23][17] ), .S(\SUMB[23][17] ) );
  FADDX1 S4_18 ( .A(\ab[23][18] ), .B(\CARRYB[22][18] ), .CI(\SUMB[22][19] ), 
        .CO(\CARRYB[23][18] ), .S(\SUMB[23][18] ) );
  FADDX1 S4_19 ( .A(\ab[23][19] ), .B(\CARRYB[22][19] ), .CI(\SUMB[22][20] ), 
        .CO(\CARRYB[23][19] ), .S(\SUMB[23][19] ) );
  FADDX1 S4_20 ( .A(\ab[23][20] ), .B(\CARRYB[22][20] ), .CI(\SUMB[22][21] ), 
        .CO(\CARRYB[23][20] ), .S(\SUMB[23][20] ) );
  FADDX1 S4_21 ( .A(\ab[23][21] ), .B(\CARRYB[22][21] ), .CI(\SUMB[22][22] ), 
        .CO(\CARRYB[23][21] ), .S(\SUMB[23][21] ) );
  FADDX1 S5_22 ( .A(\ab[23][22] ), .B(\CARRYB[22][22] ), .CI(\ab[22][23] ), 
        .CO(\CARRYB[23][22] ), .S(\SUMB[23][22] ) );
  FADDX1 S1_22_0 ( .A(\ab[22][0] ), .B(\CARRYB[21][0] ), .CI(\SUMB[21][1] ), 
        .CO(\CARRYB[22][0] ), .S(\A1[20] ) );
  FADDX1 S2_22_1 ( .A(\ab[22][1] ), .B(\CARRYB[21][1] ), .CI(\SUMB[21][2] ), 
        .CO(\CARRYB[22][1] ), .S(\SUMB[22][1] ) );
  FADDX1 S2_22_2 ( .A(\ab[22][2] ), .B(\CARRYB[21][2] ), .CI(\SUMB[21][3] ), 
        .CO(\CARRYB[22][2] ), .S(\SUMB[22][2] ) );
  FADDX1 S2_22_3 ( .A(\ab[22][3] ), .B(\CARRYB[21][3] ), .CI(\SUMB[21][4] ), 
        .CO(\CARRYB[22][3] ), .S(\SUMB[22][3] ) );
  FADDX1 S2_22_4 ( .A(\ab[22][4] ), .B(\CARRYB[21][4] ), .CI(\SUMB[21][5] ), 
        .CO(\CARRYB[22][4] ), .S(\SUMB[22][4] ) );
  FADDX1 S2_22_5 ( .A(\ab[22][5] ), .B(\CARRYB[21][5] ), .CI(\SUMB[21][6] ), 
        .CO(\CARRYB[22][5] ), .S(\SUMB[22][5] ) );
  FADDX1 S2_22_6 ( .A(\ab[22][6] ), .B(\CARRYB[21][6] ), .CI(\SUMB[21][7] ), 
        .CO(\CARRYB[22][6] ), .S(\SUMB[22][6] ) );
  FADDX1 S2_22_7 ( .A(\ab[22][7] ), .B(\CARRYB[21][7] ), .CI(\SUMB[21][8] ), 
        .CO(\CARRYB[22][7] ), .S(\SUMB[22][7] ) );
  FADDX1 S2_22_8 ( .A(\ab[22][8] ), .B(\CARRYB[21][8] ), .CI(\SUMB[21][9] ), 
        .CO(\CARRYB[22][8] ), .S(\SUMB[22][8] ) );
  FADDX1 S2_22_9 ( .A(\ab[22][9] ), .B(\CARRYB[21][9] ), .CI(\SUMB[21][10] ), 
        .CO(\CARRYB[22][9] ), .S(\SUMB[22][9] ) );
  FADDX1 S2_22_10 ( .A(\ab[22][10] ), .B(\CARRYB[21][10] ), .CI(\SUMB[21][11] ), .CO(\CARRYB[22][10] ), .S(\SUMB[22][10] ) );
  FADDX1 S2_22_11 ( .A(\ab[22][11] ), .B(\CARRYB[21][11] ), .CI(\SUMB[21][12] ), .CO(\CARRYB[22][11] ), .S(\SUMB[22][11] ) );
  FADDX1 S2_22_12 ( .A(\ab[22][12] ), .B(\CARRYB[21][12] ), .CI(\SUMB[21][13] ), .CO(\CARRYB[22][12] ), .S(\SUMB[22][12] ) );
  FADDX1 S2_22_13 ( .A(\ab[22][13] ), .B(\CARRYB[21][13] ), .CI(\SUMB[21][14] ), .CO(\CARRYB[22][13] ), .S(\SUMB[22][13] ) );
  FADDX1 S2_22_14 ( .A(\ab[22][14] ), .B(\CARRYB[21][14] ), .CI(\SUMB[21][15] ), .CO(\CARRYB[22][14] ), .S(\SUMB[22][14] ) );
  FADDX1 S2_22_15 ( .A(\ab[22][15] ), .B(\CARRYB[21][15] ), .CI(\SUMB[21][16] ), .CO(\CARRYB[22][15] ), .S(\SUMB[22][15] ) );
  FADDX1 S2_22_16 ( .A(\ab[22][16] ), .B(\CARRYB[21][16] ), .CI(\SUMB[21][17] ), .CO(\CARRYB[22][16] ), .S(\SUMB[22][16] ) );
  FADDX1 S2_22_17 ( .A(\ab[22][17] ), .B(\CARRYB[21][17] ), .CI(\SUMB[21][18] ), .CO(\CARRYB[22][17] ), .S(\SUMB[22][17] ) );
  FADDX1 S2_22_18 ( .A(\ab[22][18] ), .B(\CARRYB[21][18] ), .CI(\SUMB[21][19] ), .CO(\CARRYB[22][18] ), .S(\SUMB[22][18] ) );
  FADDX1 S2_22_19 ( .A(\ab[22][19] ), .B(\CARRYB[21][19] ), .CI(\SUMB[21][20] ), .CO(\CARRYB[22][19] ), .S(\SUMB[22][19] ) );
  FADDX1 S2_22_20 ( .A(\ab[22][20] ), .B(\CARRYB[21][20] ), .CI(\SUMB[21][21] ), .CO(\CARRYB[22][20] ), .S(\SUMB[22][20] ) );
  FADDX1 S2_22_21 ( .A(\ab[22][21] ), .B(\CARRYB[21][21] ), .CI(\SUMB[21][22] ), .CO(\CARRYB[22][21] ), .S(\SUMB[22][21] ) );
  FADDX1 S3_22_22 ( .A(\ab[22][22] ), .B(\CARRYB[21][22] ), .CI(\ab[21][23] ), 
        .CO(\CARRYB[22][22] ), .S(\SUMB[22][22] ) );
  FADDX1 S1_21_0 ( .A(\ab[21][0] ), .B(\CARRYB[20][0] ), .CI(\SUMB[20][1] ), 
        .CO(\CARRYB[21][0] ), .S(\A1[19] ) );
  FADDX1 S2_21_1 ( .A(\ab[21][1] ), .B(\CARRYB[20][1] ), .CI(\SUMB[20][2] ), 
        .CO(\CARRYB[21][1] ), .S(\SUMB[21][1] ) );
  FADDX1 S2_21_2 ( .A(\ab[21][2] ), .B(\CARRYB[20][2] ), .CI(\SUMB[20][3] ), 
        .CO(\CARRYB[21][2] ), .S(\SUMB[21][2] ) );
  FADDX1 S2_21_3 ( .A(\ab[21][3] ), .B(\CARRYB[20][3] ), .CI(\SUMB[20][4] ), 
        .CO(\CARRYB[21][3] ), .S(\SUMB[21][3] ) );
  FADDX1 S2_21_4 ( .A(\ab[21][4] ), .B(\CARRYB[20][4] ), .CI(\SUMB[20][5] ), 
        .CO(\CARRYB[21][4] ), .S(\SUMB[21][4] ) );
  FADDX1 S2_21_5 ( .A(\ab[21][5] ), .B(\CARRYB[20][5] ), .CI(\SUMB[20][6] ), 
        .CO(\CARRYB[21][5] ), .S(\SUMB[21][5] ) );
  FADDX1 S2_21_6 ( .A(\ab[21][6] ), .B(\CARRYB[20][6] ), .CI(\SUMB[20][7] ), 
        .CO(\CARRYB[21][6] ), .S(\SUMB[21][6] ) );
  FADDX1 S2_21_7 ( .A(\ab[21][7] ), .B(\CARRYB[20][7] ), .CI(\SUMB[20][8] ), 
        .CO(\CARRYB[21][7] ), .S(\SUMB[21][7] ) );
  FADDX1 S2_21_8 ( .A(\ab[21][8] ), .B(\CARRYB[20][8] ), .CI(\SUMB[20][9] ), 
        .CO(\CARRYB[21][8] ), .S(\SUMB[21][8] ) );
  FADDX1 S2_21_9 ( .A(\ab[21][9] ), .B(\CARRYB[20][9] ), .CI(\SUMB[20][10] ), 
        .CO(\CARRYB[21][9] ), .S(\SUMB[21][9] ) );
  FADDX1 S2_21_10 ( .A(\ab[21][10] ), .B(\CARRYB[20][10] ), .CI(\SUMB[20][11] ), .CO(\CARRYB[21][10] ), .S(\SUMB[21][10] ) );
  FADDX1 S2_21_11 ( .A(\ab[21][11] ), .B(\CARRYB[20][11] ), .CI(\SUMB[20][12] ), .CO(\CARRYB[21][11] ), .S(\SUMB[21][11] ) );
  FADDX1 S2_21_12 ( .A(\ab[21][12] ), .B(\CARRYB[20][12] ), .CI(\SUMB[20][13] ), .CO(\CARRYB[21][12] ), .S(\SUMB[21][12] ) );
  FADDX1 S2_21_13 ( .A(\ab[21][13] ), .B(\CARRYB[20][13] ), .CI(\SUMB[20][14] ), .CO(\CARRYB[21][13] ), .S(\SUMB[21][13] ) );
  FADDX1 S2_21_14 ( .A(\ab[21][14] ), .B(\CARRYB[20][14] ), .CI(\SUMB[20][15] ), .CO(\CARRYB[21][14] ), .S(\SUMB[21][14] ) );
  FADDX1 S2_21_15 ( .A(\ab[21][15] ), .B(\CARRYB[20][15] ), .CI(\SUMB[20][16] ), .CO(\CARRYB[21][15] ), .S(\SUMB[21][15] ) );
  FADDX1 S2_21_16 ( .A(\ab[21][16] ), .B(\CARRYB[20][16] ), .CI(\SUMB[20][17] ), .CO(\CARRYB[21][16] ), .S(\SUMB[21][16] ) );
  FADDX1 S2_21_17 ( .A(\ab[21][17] ), .B(\CARRYB[20][17] ), .CI(\SUMB[20][18] ), .CO(\CARRYB[21][17] ), .S(\SUMB[21][17] ) );
  FADDX1 S2_21_18 ( .A(\ab[21][18] ), .B(\CARRYB[20][18] ), .CI(\SUMB[20][19] ), .CO(\CARRYB[21][18] ), .S(\SUMB[21][18] ) );
  FADDX1 S2_21_19 ( .A(\ab[21][19] ), .B(\CARRYB[20][19] ), .CI(\SUMB[20][20] ), .CO(\CARRYB[21][19] ), .S(\SUMB[21][19] ) );
  FADDX1 S2_21_20 ( .A(\ab[21][20] ), .B(\CARRYB[20][20] ), .CI(\SUMB[20][21] ), .CO(\CARRYB[21][20] ), .S(\SUMB[21][20] ) );
  FADDX1 S2_21_21 ( .A(\ab[21][21] ), .B(\CARRYB[20][21] ), .CI(\SUMB[20][22] ), .CO(\CARRYB[21][21] ), .S(\SUMB[21][21] ) );
  FADDX1 S3_21_22 ( .A(\ab[21][22] ), .B(\CARRYB[20][22] ), .CI(\ab[20][23] ), 
        .CO(\CARRYB[21][22] ), .S(\SUMB[21][22] ) );
  FADDX1 S1_20_0 ( .A(\ab[20][0] ), .B(\CARRYB[19][0] ), .CI(\SUMB[19][1] ), 
        .CO(\CARRYB[20][0] ), .S(\A1[18] ) );
  FADDX1 S2_20_1 ( .A(\ab[20][1] ), .B(\CARRYB[19][1] ), .CI(\SUMB[19][2] ), 
        .CO(\CARRYB[20][1] ), .S(\SUMB[20][1] ) );
  FADDX1 S2_20_2 ( .A(\ab[20][2] ), .B(\CARRYB[19][2] ), .CI(\SUMB[19][3] ), 
        .CO(\CARRYB[20][2] ), .S(\SUMB[20][2] ) );
  FADDX1 S2_20_3 ( .A(\ab[20][3] ), .B(\CARRYB[19][3] ), .CI(\SUMB[19][4] ), 
        .CO(\CARRYB[20][3] ), .S(\SUMB[20][3] ) );
  FADDX1 S2_20_4 ( .A(\ab[20][4] ), .B(\CARRYB[19][4] ), .CI(\SUMB[19][5] ), 
        .CO(\CARRYB[20][4] ), .S(\SUMB[20][4] ) );
  FADDX1 S2_20_5 ( .A(\ab[20][5] ), .B(\CARRYB[19][5] ), .CI(\SUMB[19][6] ), 
        .CO(\CARRYB[20][5] ), .S(\SUMB[20][5] ) );
  FADDX1 S2_20_6 ( .A(\ab[20][6] ), .B(\CARRYB[19][6] ), .CI(\SUMB[19][7] ), 
        .CO(\CARRYB[20][6] ), .S(\SUMB[20][6] ) );
  FADDX1 S2_20_7 ( .A(\ab[20][7] ), .B(\CARRYB[19][7] ), .CI(\SUMB[19][8] ), 
        .CO(\CARRYB[20][7] ), .S(\SUMB[20][7] ) );
  FADDX1 S2_20_8 ( .A(\ab[20][8] ), .B(\CARRYB[19][8] ), .CI(\SUMB[19][9] ), 
        .CO(\CARRYB[20][8] ), .S(\SUMB[20][8] ) );
  FADDX1 S2_20_9 ( .A(\ab[20][9] ), .B(\CARRYB[19][9] ), .CI(\SUMB[19][10] ), 
        .CO(\CARRYB[20][9] ), .S(\SUMB[20][9] ) );
  FADDX1 S2_20_10 ( .A(\ab[20][10] ), .B(\CARRYB[19][10] ), .CI(\SUMB[19][11] ), .CO(\CARRYB[20][10] ), .S(\SUMB[20][10] ) );
  FADDX1 S2_20_11 ( .A(\ab[20][11] ), .B(\CARRYB[19][11] ), .CI(\SUMB[19][12] ), .CO(\CARRYB[20][11] ), .S(\SUMB[20][11] ) );
  FADDX1 S2_20_12 ( .A(\ab[20][12] ), .B(\CARRYB[19][12] ), .CI(\SUMB[19][13] ), .CO(\CARRYB[20][12] ), .S(\SUMB[20][12] ) );
  FADDX1 S2_20_13 ( .A(\ab[20][13] ), .B(\CARRYB[19][13] ), .CI(\SUMB[19][14] ), .CO(\CARRYB[20][13] ), .S(\SUMB[20][13] ) );
  FADDX1 S2_20_14 ( .A(\ab[20][14] ), .B(\CARRYB[19][14] ), .CI(\SUMB[19][15] ), .CO(\CARRYB[20][14] ), .S(\SUMB[20][14] ) );
  FADDX1 S2_20_15 ( .A(\ab[20][15] ), .B(\CARRYB[19][15] ), .CI(\SUMB[19][16] ), .CO(\CARRYB[20][15] ), .S(\SUMB[20][15] ) );
  FADDX1 S2_20_16 ( .A(\ab[20][16] ), .B(\CARRYB[19][16] ), .CI(\SUMB[19][17] ), .CO(\CARRYB[20][16] ), .S(\SUMB[20][16] ) );
  FADDX1 S2_20_17 ( .A(\ab[20][17] ), .B(\CARRYB[19][17] ), .CI(\SUMB[19][18] ), .CO(\CARRYB[20][17] ), .S(\SUMB[20][17] ) );
  FADDX1 S2_20_18 ( .A(\ab[20][18] ), .B(\CARRYB[19][18] ), .CI(\SUMB[19][19] ), .CO(\CARRYB[20][18] ), .S(\SUMB[20][18] ) );
  FADDX1 S2_20_19 ( .A(\ab[20][19] ), .B(\CARRYB[19][19] ), .CI(\SUMB[19][20] ), .CO(\CARRYB[20][19] ), .S(\SUMB[20][19] ) );
  FADDX1 S2_20_20 ( .A(\ab[20][20] ), .B(\CARRYB[19][20] ), .CI(\SUMB[19][21] ), .CO(\CARRYB[20][20] ), .S(\SUMB[20][20] ) );
  FADDX1 S2_20_21 ( .A(\ab[20][21] ), .B(\CARRYB[19][21] ), .CI(\SUMB[19][22] ), .CO(\CARRYB[20][21] ), .S(\SUMB[20][21] ) );
  FADDX1 S3_20_22 ( .A(\ab[20][22] ), .B(\CARRYB[19][22] ), .CI(\ab[19][23] ), 
        .CO(\CARRYB[20][22] ), .S(\SUMB[20][22] ) );
  FADDX1 S1_19_0 ( .A(\ab[19][0] ), .B(\CARRYB[18][0] ), .CI(\SUMB[18][1] ), 
        .CO(\CARRYB[19][0] ), .S(\A1[17] ) );
  FADDX1 S2_19_1 ( .A(\ab[19][1] ), .B(\CARRYB[18][1] ), .CI(\SUMB[18][2] ), 
        .CO(\CARRYB[19][1] ), .S(\SUMB[19][1] ) );
  FADDX1 S2_19_2 ( .A(\ab[19][2] ), .B(\CARRYB[18][2] ), .CI(\SUMB[18][3] ), 
        .CO(\CARRYB[19][2] ), .S(\SUMB[19][2] ) );
  FADDX1 S2_19_3 ( .A(\ab[19][3] ), .B(\CARRYB[18][3] ), .CI(\SUMB[18][4] ), 
        .CO(\CARRYB[19][3] ), .S(\SUMB[19][3] ) );
  FADDX1 S2_19_4 ( .A(\ab[19][4] ), .B(\CARRYB[18][4] ), .CI(\SUMB[18][5] ), 
        .CO(\CARRYB[19][4] ), .S(\SUMB[19][4] ) );
  FADDX1 S2_19_5 ( .A(\ab[19][5] ), .B(\CARRYB[18][5] ), .CI(\SUMB[18][6] ), 
        .CO(\CARRYB[19][5] ), .S(\SUMB[19][5] ) );
  FADDX1 S2_19_6 ( .A(\ab[19][6] ), .B(\CARRYB[18][6] ), .CI(\SUMB[18][7] ), 
        .CO(\CARRYB[19][6] ), .S(\SUMB[19][6] ) );
  FADDX1 S2_19_7 ( .A(\ab[19][7] ), .B(\CARRYB[18][7] ), .CI(\SUMB[18][8] ), 
        .CO(\CARRYB[19][7] ), .S(\SUMB[19][7] ) );
  FADDX1 S2_19_8 ( .A(\ab[19][8] ), .B(\CARRYB[18][8] ), .CI(\SUMB[18][9] ), 
        .CO(\CARRYB[19][8] ), .S(\SUMB[19][8] ) );
  FADDX1 S2_19_9 ( .A(\ab[19][9] ), .B(\CARRYB[18][9] ), .CI(\SUMB[18][10] ), 
        .CO(\CARRYB[19][9] ), .S(\SUMB[19][9] ) );
  FADDX1 S2_19_10 ( .A(\ab[19][10] ), .B(\CARRYB[18][10] ), .CI(\SUMB[18][11] ), .CO(\CARRYB[19][10] ), .S(\SUMB[19][10] ) );
  FADDX1 S2_19_11 ( .A(\ab[19][11] ), .B(\CARRYB[18][11] ), .CI(\SUMB[18][12] ), .CO(\CARRYB[19][11] ), .S(\SUMB[19][11] ) );
  FADDX1 S2_19_12 ( .A(\ab[19][12] ), .B(\CARRYB[18][12] ), .CI(\SUMB[18][13] ), .CO(\CARRYB[19][12] ), .S(\SUMB[19][12] ) );
  FADDX1 S2_19_13 ( .A(\ab[19][13] ), .B(\CARRYB[18][13] ), .CI(\SUMB[18][14] ), .CO(\CARRYB[19][13] ), .S(\SUMB[19][13] ) );
  FADDX1 S2_19_14 ( .A(\ab[19][14] ), .B(\CARRYB[18][14] ), .CI(\SUMB[18][15] ), .CO(\CARRYB[19][14] ), .S(\SUMB[19][14] ) );
  FADDX1 S2_19_15 ( .A(\ab[19][15] ), .B(\CARRYB[18][15] ), .CI(\SUMB[18][16] ), .CO(\CARRYB[19][15] ), .S(\SUMB[19][15] ) );
  FADDX1 S2_19_16 ( .A(\ab[19][16] ), .B(\CARRYB[18][16] ), .CI(\SUMB[18][17] ), .CO(\CARRYB[19][16] ), .S(\SUMB[19][16] ) );
  FADDX1 S2_19_17 ( .A(\ab[19][17] ), .B(\CARRYB[18][17] ), .CI(\SUMB[18][18] ), .CO(\CARRYB[19][17] ), .S(\SUMB[19][17] ) );
  FADDX1 S2_19_18 ( .A(\ab[19][18] ), .B(\CARRYB[18][18] ), .CI(\SUMB[18][19] ), .CO(\CARRYB[19][18] ), .S(\SUMB[19][18] ) );
  FADDX1 S2_19_19 ( .A(\ab[19][19] ), .B(\CARRYB[18][19] ), .CI(\SUMB[18][20] ), .CO(\CARRYB[19][19] ), .S(\SUMB[19][19] ) );
  FADDX1 S2_19_20 ( .A(\ab[19][20] ), .B(\CARRYB[18][20] ), .CI(\SUMB[18][21] ), .CO(\CARRYB[19][20] ), .S(\SUMB[19][20] ) );
  FADDX1 S2_19_21 ( .A(\ab[19][21] ), .B(\CARRYB[18][21] ), .CI(\SUMB[18][22] ), .CO(\CARRYB[19][21] ), .S(\SUMB[19][21] ) );
  FADDX1 S3_19_22 ( .A(\ab[19][22] ), .B(\CARRYB[18][22] ), .CI(\ab[18][23] ), 
        .CO(\CARRYB[19][22] ), .S(\SUMB[19][22] ) );
  FADDX1 S1_18_0 ( .A(\ab[18][0] ), .B(\CARRYB[17][0] ), .CI(\SUMB[17][1] ), 
        .CO(\CARRYB[18][0] ), .S(\A1[16] ) );
  FADDX1 S2_18_1 ( .A(\ab[18][1] ), .B(\CARRYB[17][1] ), .CI(\SUMB[17][2] ), 
        .CO(\CARRYB[18][1] ), .S(\SUMB[18][1] ) );
  FADDX1 S2_18_2 ( .A(\ab[18][2] ), .B(\CARRYB[17][2] ), .CI(\SUMB[17][3] ), 
        .CO(\CARRYB[18][2] ), .S(\SUMB[18][2] ) );
  FADDX1 S2_18_3 ( .A(\ab[18][3] ), .B(\CARRYB[17][3] ), .CI(\SUMB[17][4] ), 
        .CO(\CARRYB[18][3] ), .S(\SUMB[18][3] ) );
  FADDX1 S2_18_4 ( .A(\ab[18][4] ), .B(\CARRYB[17][4] ), .CI(\SUMB[17][5] ), 
        .CO(\CARRYB[18][4] ), .S(\SUMB[18][4] ) );
  FADDX1 S2_18_5 ( .A(\ab[18][5] ), .B(\CARRYB[17][5] ), .CI(\SUMB[17][6] ), 
        .CO(\CARRYB[18][5] ), .S(\SUMB[18][5] ) );
  FADDX1 S2_18_6 ( .A(\ab[18][6] ), .B(\CARRYB[17][6] ), .CI(\SUMB[17][7] ), 
        .CO(\CARRYB[18][6] ), .S(\SUMB[18][6] ) );
  FADDX1 S2_18_7 ( .A(\ab[18][7] ), .B(\CARRYB[17][7] ), .CI(\SUMB[17][8] ), 
        .CO(\CARRYB[18][7] ), .S(\SUMB[18][7] ) );
  FADDX1 S2_18_8 ( .A(\ab[18][8] ), .B(\CARRYB[17][8] ), .CI(\SUMB[17][9] ), 
        .CO(\CARRYB[18][8] ), .S(\SUMB[18][8] ) );
  FADDX1 S2_18_9 ( .A(\ab[18][9] ), .B(\CARRYB[17][9] ), .CI(\SUMB[17][10] ), 
        .CO(\CARRYB[18][9] ), .S(\SUMB[18][9] ) );
  FADDX1 S2_18_10 ( .A(\ab[18][10] ), .B(\CARRYB[17][10] ), .CI(\SUMB[17][11] ), .CO(\CARRYB[18][10] ), .S(\SUMB[18][10] ) );
  FADDX1 S2_18_11 ( .A(\ab[18][11] ), .B(\CARRYB[17][11] ), .CI(\SUMB[17][12] ), .CO(\CARRYB[18][11] ), .S(\SUMB[18][11] ) );
  FADDX1 S2_18_12 ( .A(\ab[18][12] ), .B(\CARRYB[17][12] ), .CI(\SUMB[17][13] ), .CO(\CARRYB[18][12] ), .S(\SUMB[18][12] ) );
  FADDX1 S2_18_13 ( .A(\ab[18][13] ), .B(\CARRYB[17][13] ), .CI(\SUMB[17][14] ), .CO(\CARRYB[18][13] ), .S(\SUMB[18][13] ) );
  FADDX1 S2_18_14 ( .A(\ab[18][14] ), .B(\CARRYB[17][14] ), .CI(\SUMB[17][15] ), .CO(\CARRYB[18][14] ), .S(\SUMB[18][14] ) );
  FADDX1 S2_18_15 ( .A(\ab[18][15] ), .B(\CARRYB[17][15] ), .CI(\SUMB[17][16] ), .CO(\CARRYB[18][15] ), .S(\SUMB[18][15] ) );
  FADDX1 S2_18_16 ( .A(\ab[18][16] ), .B(\CARRYB[17][16] ), .CI(\SUMB[17][17] ), .CO(\CARRYB[18][16] ), .S(\SUMB[18][16] ) );
  FADDX1 S2_18_17 ( .A(\ab[18][17] ), .B(\CARRYB[17][17] ), .CI(\SUMB[17][18] ), .CO(\CARRYB[18][17] ), .S(\SUMB[18][17] ) );
  FADDX1 S2_18_18 ( .A(\ab[18][18] ), .B(\CARRYB[17][18] ), .CI(\SUMB[17][19] ), .CO(\CARRYB[18][18] ), .S(\SUMB[18][18] ) );
  FADDX1 S2_18_19 ( .A(\ab[18][19] ), .B(\CARRYB[17][19] ), .CI(\SUMB[17][20] ), .CO(\CARRYB[18][19] ), .S(\SUMB[18][19] ) );
  FADDX1 S2_18_20 ( .A(\ab[18][20] ), .B(\CARRYB[17][20] ), .CI(\SUMB[17][21] ), .CO(\CARRYB[18][20] ), .S(\SUMB[18][20] ) );
  FADDX1 S2_18_21 ( .A(\ab[18][21] ), .B(\CARRYB[17][21] ), .CI(\SUMB[17][22] ), .CO(\CARRYB[18][21] ), .S(\SUMB[18][21] ) );
  FADDX1 S3_18_22 ( .A(\ab[18][22] ), .B(\CARRYB[17][22] ), .CI(\ab[17][23] ), 
        .CO(\CARRYB[18][22] ), .S(\SUMB[18][22] ) );
  FADDX1 S1_17_0 ( .A(\ab[17][0] ), .B(\CARRYB[16][0] ), .CI(\SUMB[16][1] ), 
        .CO(\CARRYB[17][0] ), .S(\A1[15] ) );
  FADDX1 S2_17_1 ( .A(\ab[17][1] ), .B(\CARRYB[16][1] ), .CI(\SUMB[16][2] ), 
        .CO(\CARRYB[17][1] ), .S(\SUMB[17][1] ) );
  FADDX1 S2_17_2 ( .A(\ab[17][2] ), .B(\CARRYB[16][2] ), .CI(\SUMB[16][3] ), 
        .CO(\CARRYB[17][2] ), .S(\SUMB[17][2] ) );
  FADDX1 S2_17_3 ( .A(\ab[17][3] ), .B(\CARRYB[16][3] ), .CI(\SUMB[16][4] ), 
        .CO(\CARRYB[17][3] ), .S(\SUMB[17][3] ) );
  FADDX1 S2_17_4 ( .A(\ab[17][4] ), .B(\CARRYB[16][4] ), .CI(\SUMB[16][5] ), 
        .CO(\CARRYB[17][4] ), .S(\SUMB[17][4] ) );
  FADDX1 S2_17_5 ( .A(\ab[17][5] ), .B(\CARRYB[16][5] ), .CI(\SUMB[16][6] ), 
        .CO(\CARRYB[17][5] ), .S(\SUMB[17][5] ) );
  FADDX1 S2_17_6 ( .A(\ab[17][6] ), .B(\CARRYB[16][6] ), .CI(\SUMB[16][7] ), 
        .CO(\CARRYB[17][6] ), .S(\SUMB[17][6] ) );
  FADDX1 S2_17_7 ( .A(\ab[17][7] ), .B(\CARRYB[16][7] ), .CI(\SUMB[16][8] ), 
        .CO(\CARRYB[17][7] ), .S(\SUMB[17][7] ) );
  FADDX1 S2_17_8 ( .A(\ab[17][8] ), .B(\CARRYB[16][8] ), .CI(\SUMB[16][9] ), 
        .CO(\CARRYB[17][8] ), .S(\SUMB[17][8] ) );
  FADDX1 S2_17_9 ( .A(\ab[17][9] ), .B(\CARRYB[16][9] ), .CI(\SUMB[16][10] ), 
        .CO(\CARRYB[17][9] ), .S(\SUMB[17][9] ) );
  FADDX1 S2_17_10 ( .A(\ab[17][10] ), .B(\CARRYB[16][10] ), .CI(\SUMB[16][11] ), .CO(\CARRYB[17][10] ), .S(\SUMB[17][10] ) );
  FADDX1 S2_17_11 ( .A(\ab[17][11] ), .B(\CARRYB[16][11] ), .CI(\SUMB[16][12] ), .CO(\CARRYB[17][11] ), .S(\SUMB[17][11] ) );
  FADDX1 S2_17_12 ( .A(\ab[17][12] ), .B(\CARRYB[16][12] ), .CI(\SUMB[16][13] ), .CO(\CARRYB[17][12] ), .S(\SUMB[17][12] ) );
  FADDX1 S2_17_13 ( .A(\ab[17][13] ), .B(\CARRYB[16][13] ), .CI(\SUMB[16][14] ), .CO(\CARRYB[17][13] ), .S(\SUMB[17][13] ) );
  FADDX1 S2_17_14 ( .A(\ab[17][14] ), .B(\CARRYB[16][14] ), .CI(\SUMB[16][15] ), .CO(\CARRYB[17][14] ), .S(\SUMB[17][14] ) );
  FADDX1 S2_17_15 ( .A(\ab[17][15] ), .B(\CARRYB[16][15] ), .CI(\SUMB[16][16] ), .CO(\CARRYB[17][15] ), .S(\SUMB[17][15] ) );
  FADDX1 S2_17_16 ( .A(\ab[17][16] ), .B(\CARRYB[16][16] ), .CI(\SUMB[16][17] ), .CO(\CARRYB[17][16] ), .S(\SUMB[17][16] ) );
  FADDX1 S2_17_17 ( .A(\ab[17][17] ), .B(\CARRYB[16][17] ), .CI(\SUMB[16][18] ), .CO(\CARRYB[17][17] ), .S(\SUMB[17][17] ) );
  FADDX1 S2_17_18 ( .A(\ab[17][18] ), .B(\CARRYB[16][18] ), .CI(\SUMB[16][19] ), .CO(\CARRYB[17][18] ), .S(\SUMB[17][18] ) );
  FADDX1 S2_17_19 ( .A(\ab[17][19] ), .B(\CARRYB[16][19] ), .CI(\SUMB[16][20] ), .CO(\CARRYB[17][19] ), .S(\SUMB[17][19] ) );
  FADDX1 S2_17_20 ( .A(\ab[17][20] ), .B(\CARRYB[16][20] ), .CI(\SUMB[16][21] ), .CO(\CARRYB[17][20] ), .S(\SUMB[17][20] ) );
  FADDX1 S2_17_21 ( .A(\ab[17][21] ), .B(\CARRYB[16][21] ), .CI(\SUMB[16][22] ), .CO(\CARRYB[17][21] ), .S(\SUMB[17][21] ) );
  FADDX1 S3_17_22 ( .A(\ab[17][22] ), .B(\CARRYB[16][22] ), .CI(\ab[16][23] ), 
        .CO(\CARRYB[17][22] ), .S(\SUMB[17][22] ) );
  FADDX1 S1_16_0 ( .A(\ab[16][0] ), .B(\CARRYB[15][0] ), .CI(\SUMB[15][1] ), 
        .CO(\CARRYB[16][0] ), .S(\A1[14] ) );
  FADDX1 S2_16_1 ( .A(\ab[16][1] ), .B(\CARRYB[15][1] ), .CI(\SUMB[15][2] ), 
        .CO(\CARRYB[16][1] ), .S(\SUMB[16][1] ) );
  FADDX1 S2_16_2 ( .A(\ab[16][2] ), .B(\CARRYB[15][2] ), .CI(\SUMB[15][3] ), 
        .CO(\CARRYB[16][2] ), .S(\SUMB[16][2] ) );
  FADDX1 S2_16_3 ( .A(\ab[16][3] ), .B(\CARRYB[15][3] ), .CI(\SUMB[15][4] ), 
        .CO(\CARRYB[16][3] ), .S(\SUMB[16][3] ) );
  FADDX1 S2_16_4 ( .A(\ab[16][4] ), .B(\CARRYB[15][4] ), .CI(\SUMB[15][5] ), 
        .CO(\CARRYB[16][4] ), .S(\SUMB[16][4] ) );
  FADDX1 S2_16_5 ( .A(\ab[16][5] ), .B(\CARRYB[15][5] ), .CI(\SUMB[15][6] ), 
        .CO(\CARRYB[16][5] ), .S(\SUMB[16][5] ) );
  FADDX1 S2_16_6 ( .A(\ab[16][6] ), .B(\CARRYB[15][6] ), .CI(\SUMB[15][7] ), 
        .CO(\CARRYB[16][6] ), .S(\SUMB[16][6] ) );
  FADDX1 S2_16_7 ( .A(\ab[16][7] ), .B(\CARRYB[15][7] ), .CI(\SUMB[15][8] ), 
        .CO(\CARRYB[16][7] ), .S(\SUMB[16][7] ) );
  FADDX1 S2_16_8 ( .A(\ab[16][8] ), .B(\CARRYB[15][8] ), .CI(\SUMB[15][9] ), 
        .CO(\CARRYB[16][8] ), .S(\SUMB[16][8] ) );
  FADDX1 S2_16_9 ( .A(\ab[16][9] ), .B(\CARRYB[15][9] ), .CI(\SUMB[15][10] ), 
        .CO(\CARRYB[16][9] ), .S(\SUMB[16][9] ) );
  FADDX1 S2_16_10 ( .A(\ab[16][10] ), .B(\CARRYB[15][10] ), .CI(\SUMB[15][11] ), .CO(\CARRYB[16][10] ), .S(\SUMB[16][10] ) );
  FADDX1 S2_16_11 ( .A(\ab[16][11] ), .B(\CARRYB[15][11] ), .CI(\SUMB[15][12] ), .CO(\CARRYB[16][11] ), .S(\SUMB[16][11] ) );
  FADDX1 S2_16_12 ( .A(\ab[16][12] ), .B(\CARRYB[15][12] ), .CI(\SUMB[15][13] ), .CO(\CARRYB[16][12] ), .S(\SUMB[16][12] ) );
  FADDX1 S2_16_13 ( .A(\ab[16][13] ), .B(\CARRYB[15][13] ), .CI(\SUMB[15][14] ), .CO(\CARRYB[16][13] ), .S(\SUMB[16][13] ) );
  FADDX1 S2_16_14 ( .A(\ab[16][14] ), .B(\CARRYB[15][14] ), .CI(\SUMB[15][15] ), .CO(\CARRYB[16][14] ), .S(\SUMB[16][14] ) );
  FADDX1 S2_16_15 ( .A(\ab[16][15] ), .B(\CARRYB[15][15] ), .CI(\SUMB[15][16] ), .CO(\CARRYB[16][15] ), .S(\SUMB[16][15] ) );
  FADDX1 S2_16_16 ( .A(\ab[16][16] ), .B(\CARRYB[15][16] ), .CI(\SUMB[15][17] ), .CO(\CARRYB[16][16] ), .S(\SUMB[16][16] ) );
  FADDX1 S2_16_17 ( .A(\ab[16][17] ), .B(\CARRYB[15][17] ), .CI(\SUMB[15][18] ), .CO(\CARRYB[16][17] ), .S(\SUMB[16][17] ) );
  FADDX1 S2_16_18 ( .A(\ab[16][18] ), .B(\CARRYB[15][18] ), .CI(\SUMB[15][19] ), .CO(\CARRYB[16][18] ), .S(\SUMB[16][18] ) );
  FADDX1 S2_16_19 ( .A(\ab[16][19] ), .B(\CARRYB[15][19] ), .CI(\SUMB[15][20] ), .CO(\CARRYB[16][19] ), .S(\SUMB[16][19] ) );
  FADDX1 S2_16_20 ( .A(\ab[16][20] ), .B(\CARRYB[15][20] ), .CI(\SUMB[15][21] ), .CO(\CARRYB[16][20] ), .S(\SUMB[16][20] ) );
  FADDX1 S2_16_21 ( .A(\ab[16][21] ), .B(\CARRYB[15][21] ), .CI(\SUMB[15][22] ), .CO(\CARRYB[16][21] ), .S(\SUMB[16][21] ) );
  FADDX1 S3_16_22 ( .A(\ab[16][22] ), .B(\CARRYB[15][22] ), .CI(\ab[15][23] ), 
        .CO(\CARRYB[16][22] ), .S(\SUMB[16][22] ) );
  FADDX1 S1_15_0 ( .A(\ab[15][0] ), .B(\CARRYB[14][0] ), .CI(\SUMB[14][1] ), 
        .CO(\CARRYB[15][0] ), .S(\A1[13] ) );
  FADDX1 S2_15_1 ( .A(\ab[15][1] ), .B(\CARRYB[14][1] ), .CI(\SUMB[14][2] ), 
        .CO(\CARRYB[15][1] ), .S(\SUMB[15][1] ) );
  FADDX1 S2_15_2 ( .A(\ab[15][2] ), .B(\CARRYB[14][2] ), .CI(\SUMB[14][3] ), 
        .CO(\CARRYB[15][2] ), .S(\SUMB[15][2] ) );
  FADDX1 S2_15_3 ( .A(\ab[15][3] ), .B(\CARRYB[14][3] ), .CI(\SUMB[14][4] ), 
        .CO(\CARRYB[15][3] ), .S(\SUMB[15][3] ) );
  FADDX1 S2_15_4 ( .A(\ab[15][4] ), .B(\CARRYB[14][4] ), .CI(\SUMB[14][5] ), 
        .CO(\CARRYB[15][4] ), .S(\SUMB[15][4] ) );
  FADDX1 S2_15_5 ( .A(\ab[15][5] ), .B(\CARRYB[14][5] ), .CI(\SUMB[14][6] ), 
        .CO(\CARRYB[15][5] ), .S(\SUMB[15][5] ) );
  FADDX1 S2_15_6 ( .A(\ab[15][6] ), .B(\CARRYB[14][6] ), .CI(\SUMB[14][7] ), 
        .CO(\CARRYB[15][6] ), .S(\SUMB[15][6] ) );
  FADDX1 S2_15_7 ( .A(\ab[15][7] ), .B(\CARRYB[14][7] ), .CI(\SUMB[14][8] ), 
        .CO(\CARRYB[15][7] ), .S(\SUMB[15][7] ) );
  FADDX1 S2_15_8 ( .A(\ab[15][8] ), .B(\CARRYB[14][8] ), .CI(\SUMB[14][9] ), 
        .CO(\CARRYB[15][8] ), .S(\SUMB[15][8] ) );
  FADDX1 S2_15_9 ( .A(\ab[15][9] ), .B(\CARRYB[14][9] ), .CI(\SUMB[14][10] ), 
        .CO(\CARRYB[15][9] ), .S(\SUMB[15][9] ) );
  FADDX1 S2_15_10 ( .A(\ab[15][10] ), .B(\CARRYB[14][10] ), .CI(\SUMB[14][11] ), .CO(\CARRYB[15][10] ), .S(\SUMB[15][10] ) );
  FADDX1 S2_15_11 ( .A(\ab[15][11] ), .B(\CARRYB[14][11] ), .CI(\SUMB[14][12] ), .CO(\CARRYB[15][11] ), .S(\SUMB[15][11] ) );
  FADDX1 S2_15_12 ( .A(\ab[15][12] ), .B(\CARRYB[14][12] ), .CI(\SUMB[14][13] ), .CO(\CARRYB[15][12] ), .S(\SUMB[15][12] ) );
  FADDX1 S2_15_13 ( .A(\ab[15][13] ), .B(\CARRYB[14][13] ), .CI(\SUMB[14][14] ), .CO(\CARRYB[15][13] ), .S(\SUMB[15][13] ) );
  FADDX1 S2_15_14 ( .A(\ab[15][14] ), .B(\CARRYB[14][14] ), .CI(\SUMB[14][15] ), .CO(\CARRYB[15][14] ), .S(\SUMB[15][14] ) );
  FADDX1 S2_15_15 ( .A(\ab[15][15] ), .B(\CARRYB[14][15] ), .CI(\SUMB[14][16] ), .CO(\CARRYB[15][15] ), .S(\SUMB[15][15] ) );
  FADDX1 S2_15_16 ( .A(\ab[15][16] ), .B(\CARRYB[14][16] ), .CI(\SUMB[14][17] ), .CO(\CARRYB[15][16] ), .S(\SUMB[15][16] ) );
  FADDX1 S2_15_17 ( .A(\ab[15][17] ), .B(\CARRYB[14][17] ), .CI(\SUMB[14][18] ), .CO(\CARRYB[15][17] ), .S(\SUMB[15][17] ) );
  FADDX1 S2_15_18 ( .A(\ab[15][18] ), .B(\CARRYB[14][18] ), .CI(\SUMB[14][19] ), .CO(\CARRYB[15][18] ), .S(\SUMB[15][18] ) );
  FADDX1 S2_15_19 ( .A(\ab[15][19] ), .B(\CARRYB[14][19] ), .CI(\SUMB[14][20] ), .CO(\CARRYB[15][19] ), .S(\SUMB[15][19] ) );
  FADDX1 S2_15_20 ( .A(\ab[15][20] ), .B(\CARRYB[14][20] ), .CI(\SUMB[14][21] ), .CO(\CARRYB[15][20] ), .S(\SUMB[15][20] ) );
  FADDX1 S2_15_21 ( .A(\ab[15][21] ), .B(\CARRYB[14][21] ), .CI(\SUMB[14][22] ), .CO(\CARRYB[15][21] ), .S(\SUMB[15][21] ) );
  FADDX1 S3_15_22 ( .A(\ab[15][22] ), .B(\CARRYB[14][22] ), .CI(\ab[14][23] ), 
        .CO(\CARRYB[15][22] ), .S(\SUMB[15][22] ) );
  FADDX1 S1_14_0 ( .A(\ab[14][0] ), .B(\CARRYB[13][0] ), .CI(\SUMB[13][1] ), 
        .CO(\CARRYB[14][0] ), .S(\A1[12] ) );
  FADDX1 S2_14_1 ( .A(\ab[14][1] ), .B(\CARRYB[13][1] ), .CI(\SUMB[13][2] ), 
        .CO(\CARRYB[14][1] ), .S(\SUMB[14][1] ) );
  FADDX1 S2_14_2 ( .A(\ab[14][2] ), .B(\CARRYB[13][2] ), .CI(\SUMB[13][3] ), 
        .CO(\CARRYB[14][2] ), .S(\SUMB[14][2] ) );
  FADDX1 S2_14_3 ( .A(\ab[14][3] ), .B(\CARRYB[13][3] ), .CI(\SUMB[13][4] ), 
        .CO(\CARRYB[14][3] ), .S(\SUMB[14][3] ) );
  FADDX1 S2_14_4 ( .A(\ab[14][4] ), .B(\CARRYB[13][4] ), .CI(\SUMB[13][5] ), 
        .CO(\CARRYB[14][4] ), .S(\SUMB[14][4] ) );
  FADDX1 S2_14_5 ( .A(\ab[14][5] ), .B(\CARRYB[13][5] ), .CI(\SUMB[13][6] ), 
        .CO(\CARRYB[14][5] ), .S(\SUMB[14][5] ) );
  FADDX1 S2_14_6 ( .A(\ab[14][6] ), .B(\CARRYB[13][6] ), .CI(\SUMB[13][7] ), 
        .CO(\CARRYB[14][6] ), .S(\SUMB[14][6] ) );
  FADDX1 S2_14_7 ( .A(\ab[14][7] ), .B(\CARRYB[13][7] ), .CI(\SUMB[13][8] ), 
        .CO(\CARRYB[14][7] ), .S(\SUMB[14][7] ) );
  FADDX1 S2_14_8 ( .A(\ab[14][8] ), .B(\CARRYB[13][8] ), .CI(\SUMB[13][9] ), 
        .CO(\CARRYB[14][8] ), .S(\SUMB[14][8] ) );
  FADDX1 S2_14_9 ( .A(\ab[14][9] ), .B(\CARRYB[13][9] ), .CI(\SUMB[13][10] ), 
        .CO(\CARRYB[14][9] ), .S(\SUMB[14][9] ) );
  FADDX1 S2_14_10 ( .A(\ab[14][10] ), .B(\CARRYB[13][10] ), .CI(\SUMB[13][11] ), .CO(\CARRYB[14][10] ), .S(\SUMB[14][10] ) );
  FADDX1 S2_14_11 ( .A(\ab[14][11] ), .B(\CARRYB[13][11] ), .CI(\SUMB[13][12] ), .CO(\CARRYB[14][11] ), .S(\SUMB[14][11] ) );
  FADDX1 S2_14_12 ( .A(\ab[14][12] ), .B(\CARRYB[13][12] ), .CI(\SUMB[13][13] ), .CO(\CARRYB[14][12] ), .S(\SUMB[14][12] ) );
  FADDX1 S2_14_13 ( .A(\ab[14][13] ), .B(\CARRYB[13][13] ), .CI(\SUMB[13][14] ), .CO(\CARRYB[14][13] ), .S(\SUMB[14][13] ) );
  FADDX1 S2_14_14 ( .A(\ab[14][14] ), .B(\CARRYB[13][14] ), .CI(\SUMB[13][15] ), .CO(\CARRYB[14][14] ), .S(\SUMB[14][14] ) );
  FADDX1 S2_14_15 ( .A(\ab[14][15] ), .B(\CARRYB[13][15] ), .CI(\SUMB[13][16] ), .CO(\CARRYB[14][15] ), .S(\SUMB[14][15] ) );
  FADDX1 S2_14_16 ( .A(\ab[14][16] ), .B(\CARRYB[13][16] ), .CI(\SUMB[13][17] ), .CO(\CARRYB[14][16] ), .S(\SUMB[14][16] ) );
  FADDX1 S2_14_17 ( .A(\ab[14][17] ), .B(\CARRYB[13][17] ), .CI(\SUMB[13][18] ), .CO(\CARRYB[14][17] ), .S(\SUMB[14][17] ) );
  FADDX1 S2_14_18 ( .A(\ab[14][18] ), .B(\CARRYB[13][18] ), .CI(\SUMB[13][19] ), .CO(\CARRYB[14][18] ), .S(\SUMB[14][18] ) );
  FADDX1 S2_14_19 ( .A(\ab[14][19] ), .B(\CARRYB[13][19] ), .CI(\SUMB[13][20] ), .CO(\CARRYB[14][19] ), .S(\SUMB[14][19] ) );
  FADDX1 S2_14_20 ( .A(\ab[14][20] ), .B(\CARRYB[13][20] ), .CI(\SUMB[13][21] ), .CO(\CARRYB[14][20] ), .S(\SUMB[14][20] ) );
  FADDX1 S2_14_21 ( .A(\ab[14][21] ), .B(\CARRYB[13][21] ), .CI(\SUMB[13][22] ), .CO(\CARRYB[14][21] ), .S(\SUMB[14][21] ) );
  FADDX1 S3_14_22 ( .A(\ab[14][22] ), .B(\CARRYB[13][22] ), .CI(\ab[13][23] ), 
        .CO(\CARRYB[14][22] ), .S(\SUMB[14][22] ) );
  FADDX1 S1_13_0 ( .A(\ab[13][0] ), .B(\CARRYB[12][0] ), .CI(\SUMB[12][1] ), 
        .CO(\CARRYB[13][0] ), .S(\A1[11] ) );
  FADDX1 S2_13_1 ( .A(\ab[13][1] ), .B(\CARRYB[12][1] ), .CI(\SUMB[12][2] ), 
        .CO(\CARRYB[13][1] ), .S(\SUMB[13][1] ) );
  FADDX1 S2_13_2 ( .A(\ab[13][2] ), .B(\CARRYB[12][2] ), .CI(\SUMB[12][3] ), 
        .CO(\CARRYB[13][2] ), .S(\SUMB[13][2] ) );
  FADDX1 S2_13_3 ( .A(\ab[13][3] ), .B(\CARRYB[12][3] ), .CI(\SUMB[12][4] ), 
        .CO(\CARRYB[13][3] ), .S(\SUMB[13][3] ) );
  FADDX1 S2_13_4 ( .A(\ab[13][4] ), .B(\CARRYB[12][4] ), .CI(\SUMB[12][5] ), 
        .CO(\CARRYB[13][4] ), .S(\SUMB[13][4] ) );
  FADDX1 S2_13_5 ( .A(\ab[13][5] ), .B(\CARRYB[12][5] ), .CI(\SUMB[12][6] ), 
        .CO(\CARRYB[13][5] ), .S(\SUMB[13][5] ) );
  FADDX1 S2_13_6 ( .A(\ab[13][6] ), .B(\CARRYB[12][6] ), .CI(\SUMB[12][7] ), 
        .CO(\CARRYB[13][6] ), .S(\SUMB[13][6] ) );
  FADDX1 S2_13_7 ( .A(\ab[13][7] ), .B(\CARRYB[12][7] ), .CI(\SUMB[12][8] ), 
        .CO(\CARRYB[13][7] ), .S(\SUMB[13][7] ) );
  FADDX1 S2_13_8 ( .A(\ab[13][8] ), .B(\CARRYB[12][8] ), .CI(\SUMB[12][9] ), 
        .CO(\CARRYB[13][8] ), .S(\SUMB[13][8] ) );
  FADDX1 S2_13_9 ( .A(\ab[13][9] ), .B(\CARRYB[12][9] ), .CI(\SUMB[12][10] ), 
        .CO(\CARRYB[13][9] ), .S(\SUMB[13][9] ) );
  FADDX1 S2_13_10 ( .A(\ab[13][10] ), .B(\CARRYB[12][10] ), .CI(\SUMB[12][11] ), .CO(\CARRYB[13][10] ), .S(\SUMB[13][10] ) );
  FADDX1 S2_13_11 ( .A(\ab[13][11] ), .B(\CARRYB[12][11] ), .CI(\SUMB[12][12] ), .CO(\CARRYB[13][11] ), .S(\SUMB[13][11] ) );
  FADDX1 S2_13_12 ( .A(\ab[13][12] ), .B(\CARRYB[12][12] ), .CI(\SUMB[12][13] ), .CO(\CARRYB[13][12] ), .S(\SUMB[13][12] ) );
  FADDX1 S2_13_13 ( .A(\ab[13][13] ), .B(\CARRYB[12][13] ), .CI(\SUMB[12][14] ), .CO(\CARRYB[13][13] ), .S(\SUMB[13][13] ) );
  FADDX1 S2_13_14 ( .A(\ab[13][14] ), .B(\CARRYB[12][14] ), .CI(\SUMB[12][15] ), .CO(\CARRYB[13][14] ), .S(\SUMB[13][14] ) );
  FADDX1 S2_13_15 ( .A(\ab[13][15] ), .B(\CARRYB[12][15] ), .CI(\SUMB[12][16] ), .CO(\CARRYB[13][15] ), .S(\SUMB[13][15] ) );
  FADDX1 S2_13_16 ( .A(\ab[13][16] ), .B(\CARRYB[12][16] ), .CI(\SUMB[12][17] ), .CO(\CARRYB[13][16] ), .S(\SUMB[13][16] ) );
  FADDX1 S2_13_17 ( .A(\ab[13][17] ), .B(\CARRYB[12][17] ), .CI(\SUMB[12][18] ), .CO(\CARRYB[13][17] ), .S(\SUMB[13][17] ) );
  FADDX1 S2_13_18 ( .A(\ab[13][18] ), .B(\CARRYB[12][18] ), .CI(\SUMB[12][19] ), .CO(\CARRYB[13][18] ), .S(\SUMB[13][18] ) );
  FADDX1 S2_13_19 ( .A(\ab[13][19] ), .B(\CARRYB[12][19] ), .CI(\SUMB[12][20] ), .CO(\CARRYB[13][19] ), .S(\SUMB[13][19] ) );
  FADDX1 S2_13_20 ( .A(\ab[13][20] ), .B(\CARRYB[12][20] ), .CI(\SUMB[12][21] ), .CO(\CARRYB[13][20] ), .S(\SUMB[13][20] ) );
  FADDX1 S2_13_21 ( .A(\ab[13][21] ), .B(\CARRYB[12][21] ), .CI(\SUMB[12][22] ), .CO(\CARRYB[13][21] ), .S(\SUMB[13][21] ) );
  FADDX1 S3_13_22 ( .A(\ab[13][22] ), .B(\CARRYB[12][22] ), .CI(\ab[12][23] ), 
        .CO(\CARRYB[13][22] ), .S(\SUMB[13][22] ) );
  FADDX1 S1_12_0 ( .A(\ab[12][0] ), .B(\CARRYB[11][0] ), .CI(\SUMB[11][1] ), 
        .CO(\CARRYB[12][0] ), .S(\A1[10] ) );
  FADDX1 S2_12_1 ( .A(\ab[12][1] ), .B(\CARRYB[11][1] ), .CI(\SUMB[11][2] ), 
        .CO(\CARRYB[12][1] ), .S(\SUMB[12][1] ) );
  FADDX1 S2_12_2 ( .A(\ab[12][2] ), .B(\CARRYB[11][2] ), .CI(\SUMB[11][3] ), 
        .CO(\CARRYB[12][2] ), .S(\SUMB[12][2] ) );
  FADDX1 S2_12_3 ( .A(\ab[12][3] ), .B(\CARRYB[11][3] ), .CI(\SUMB[11][4] ), 
        .CO(\CARRYB[12][3] ), .S(\SUMB[12][3] ) );
  FADDX1 S2_12_4 ( .A(\ab[12][4] ), .B(\CARRYB[11][4] ), .CI(\SUMB[11][5] ), 
        .CO(\CARRYB[12][4] ), .S(\SUMB[12][4] ) );
  FADDX1 S2_12_5 ( .A(\ab[12][5] ), .B(\CARRYB[11][5] ), .CI(\SUMB[11][6] ), 
        .CO(\CARRYB[12][5] ), .S(\SUMB[12][5] ) );
  FADDX1 S2_12_6 ( .A(\ab[12][6] ), .B(\CARRYB[11][6] ), .CI(\SUMB[11][7] ), 
        .CO(\CARRYB[12][6] ), .S(\SUMB[12][6] ) );
  FADDX1 S2_12_7 ( .A(\ab[12][7] ), .B(\CARRYB[11][7] ), .CI(\SUMB[11][8] ), 
        .CO(\CARRYB[12][7] ), .S(\SUMB[12][7] ) );
  FADDX1 S2_12_8 ( .A(\ab[12][8] ), .B(\CARRYB[11][8] ), .CI(\SUMB[11][9] ), 
        .CO(\CARRYB[12][8] ), .S(\SUMB[12][8] ) );
  FADDX1 S2_12_9 ( .A(\ab[12][9] ), .B(\CARRYB[11][9] ), .CI(\SUMB[11][10] ), 
        .CO(\CARRYB[12][9] ), .S(\SUMB[12][9] ) );
  FADDX1 S2_12_10 ( .A(\ab[12][10] ), .B(\CARRYB[11][10] ), .CI(\SUMB[11][11] ), .CO(\CARRYB[12][10] ), .S(\SUMB[12][10] ) );
  FADDX1 S2_12_11 ( .A(\ab[12][11] ), .B(\CARRYB[11][11] ), .CI(\SUMB[11][12] ), .CO(\CARRYB[12][11] ), .S(\SUMB[12][11] ) );
  FADDX1 S2_12_12 ( .A(\ab[12][12] ), .B(\CARRYB[11][12] ), .CI(\SUMB[11][13] ), .CO(\CARRYB[12][12] ), .S(\SUMB[12][12] ) );
  FADDX1 S2_12_13 ( .A(\ab[12][13] ), .B(\CARRYB[11][13] ), .CI(\SUMB[11][14] ), .CO(\CARRYB[12][13] ), .S(\SUMB[12][13] ) );
  FADDX1 S2_12_14 ( .A(\ab[12][14] ), .B(\CARRYB[11][14] ), .CI(\SUMB[11][15] ), .CO(\CARRYB[12][14] ), .S(\SUMB[12][14] ) );
  FADDX1 S2_12_15 ( .A(\ab[12][15] ), .B(\CARRYB[11][15] ), .CI(\SUMB[11][16] ), .CO(\CARRYB[12][15] ), .S(\SUMB[12][15] ) );
  FADDX1 S2_12_16 ( .A(\ab[12][16] ), .B(\CARRYB[11][16] ), .CI(\SUMB[11][17] ), .CO(\CARRYB[12][16] ), .S(\SUMB[12][16] ) );
  FADDX1 S2_12_17 ( .A(\ab[12][17] ), .B(\CARRYB[11][17] ), .CI(\SUMB[11][18] ), .CO(\CARRYB[12][17] ), .S(\SUMB[12][17] ) );
  FADDX1 S2_12_18 ( .A(\ab[12][18] ), .B(\CARRYB[11][18] ), .CI(\SUMB[11][19] ), .CO(\CARRYB[12][18] ), .S(\SUMB[12][18] ) );
  FADDX1 S2_12_19 ( .A(\ab[12][19] ), .B(\CARRYB[11][19] ), .CI(\SUMB[11][20] ), .CO(\CARRYB[12][19] ), .S(\SUMB[12][19] ) );
  FADDX1 S2_12_20 ( .A(\ab[12][20] ), .B(\CARRYB[11][20] ), .CI(\SUMB[11][21] ), .CO(\CARRYB[12][20] ), .S(\SUMB[12][20] ) );
  FADDX1 S2_12_21 ( .A(\ab[12][21] ), .B(\CARRYB[11][21] ), .CI(\SUMB[11][22] ), .CO(\CARRYB[12][21] ), .S(\SUMB[12][21] ) );
  FADDX1 S3_12_22 ( .A(\ab[12][22] ), .B(\CARRYB[11][22] ), .CI(\ab[11][23] ), 
        .CO(\CARRYB[12][22] ), .S(\SUMB[12][22] ) );
  FADDX1 S1_11_0 ( .A(\ab[11][0] ), .B(\CARRYB[10][0] ), .CI(\SUMB[10][1] ), 
        .CO(\CARRYB[11][0] ), .S(\A1[9] ) );
  FADDX1 S2_11_1 ( .A(\ab[11][1] ), .B(\CARRYB[10][1] ), .CI(\SUMB[10][2] ), 
        .CO(\CARRYB[11][1] ), .S(\SUMB[11][1] ) );
  FADDX1 S2_11_2 ( .A(\ab[11][2] ), .B(\CARRYB[10][2] ), .CI(\SUMB[10][3] ), 
        .CO(\CARRYB[11][2] ), .S(\SUMB[11][2] ) );
  FADDX1 S2_11_3 ( .A(\ab[11][3] ), .B(\CARRYB[10][3] ), .CI(\SUMB[10][4] ), 
        .CO(\CARRYB[11][3] ), .S(\SUMB[11][3] ) );
  FADDX1 S2_11_4 ( .A(\ab[11][4] ), .B(\CARRYB[10][4] ), .CI(\SUMB[10][5] ), 
        .CO(\CARRYB[11][4] ), .S(\SUMB[11][4] ) );
  FADDX1 S2_11_5 ( .A(\ab[11][5] ), .B(\CARRYB[10][5] ), .CI(\SUMB[10][6] ), 
        .CO(\CARRYB[11][5] ), .S(\SUMB[11][5] ) );
  FADDX1 S2_11_6 ( .A(\ab[11][6] ), .B(\CARRYB[10][6] ), .CI(\SUMB[10][7] ), 
        .CO(\CARRYB[11][6] ), .S(\SUMB[11][6] ) );
  FADDX1 S2_11_7 ( .A(\ab[11][7] ), .B(\CARRYB[10][7] ), .CI(\SUMB[10][8] ), 
        .CO(\CARRYB[11][7] ), .S(\SUMB[11][7] ) );
  FADDX1 S2_11_8 ( .A(\ab[11][8] ), .B(\CARRYB[10][8] ), .CI(\SUMB[10][9] ), 
        .CO(\CARRYB[11][8] ), .S(\SUMB[11][8] ) );
  FADDX1 S2_11_9 ( .A(\ab[11][9] ), .B(\CARRYB[10][9] ), .CI(\SUMB[10][10] ), 
        .CO(\CARRYB[11][9] ), .S(\SUMB[11][9] ) );
  FADDX1 S2_11_10 ( .A(\ab[11][10] ), .B(\CARRYB[10][10] ), .CI(\SUMB[10][11] ), .CO(\CARRYB[11][10] ), .S(\SUMB[11][10] ) );
  FADDX1 S2_11_11 ( .A(\ab[11][11] ), .B(\CARRYB[10][11] ), .CI(\SUMB[10][12] ), .CO(\CARRYB[11][11] ), .S(\SUMB[11][11] ) );
  FADDX1 S2_11_12 ( .A(\ab[11][12] ), .B(\CARRYB[10][12] ), .CI(\SUMB[10][13] ), .CO(\CARRYB[11][12] ), .S(\SUMB[11][12] ) );
  FADDX1 S2_11_13 ( .A(\ab[11][13] ), .B(\CARRYB[10][13] ), .CI(\SUMB[10][14] ), .CO(\CARRYB[11][13] ), .S(\SUMB[11][13] ) );
  FADDX1 S2_11_14 ( .A(\ab[11][14] ), .B(\CARRYB[10][14] ), .CI(\SUMB[10][15] ), .CO(\CARRYB[11][14] ), .S(\SUMB[11][14] ) );
  FADDX1 S2_11_15 ( .A(\ab[11][15] ), .B(\CARRYB[10][15] ), .CI(\SUMB[10][16] ), .CO(\CARRYB[11][15] ), .S(\SUMB[11][15] ) );
  FADDX1 S2_11_16 ( .A(\ab[11][16] ), .B(\CARRYB[10][16] ), .CI(\SUMB[10][17] ), .CO(\CARRYB[11][16] ), .S(\SUMB[11][16] ) );
  FADDX1 S2_11_17 ( .A(\ab[11][17] ), .B(\CARRYB[10][17] ), .CI(\SUMB[10][18] ), .CO(\CARRYB[11][17] ), .S(\SUMB[11][17] ) );
  FADDX1 S2_11_18 ( .A(\ab[11][18] ), .B(\CARRYB[10][18] ), .CI(\SUMB[10][19] ), .CO(\CARRYB[11][18] ), .S(\SUMB[11][18] ) );
  FADDX1 S2_11_19 ( .A(\ab[11][19] ), .B(\CARRYB[10][19] ), .CI(\SUMB[10][20] ), .CO(\CARRYB[11][19] ), .S(\SUMB[11][19] ) );
  FADDX1 S2_11_20 ( .A(\ab[11][20] ), .B(\CARRYB[10][20] ), .CI(\SUMB[10][21] ), .CO(\CARRYB[11][20] ), .S(\SUMB[11][20] ) );
  FADDX1 S2_11_21 ( .A(\ab[11][21] ), .B(\CARRYB[10][21] ), .CI(\SUMB[10][22] ), .CO(\CARRYB[11][21] ), .S(\SUMB[11][21] ) );
  FADDX1 S3_11_22 ( .A(\ab[11][22] ), .B(\CARRYB[10][22] ), .CI(\ab[10][23] ), 
        .CO(\CARRYB[11][22] ), .S(\SUMB[11][22] ) );
  FADDX1 S1_10_0 ( .A(\ab[10][0] ), .B(\CARRYB[9][0] ), .CI(\SUMB[9][1] ), 
        .CO(\CARRYB[10][0] ), .S(\A1[8] ) );
  FADDX1 S2_10_1 ( .A(\ab[10][1] ), .B(\CARRYB[9][1] ), .CI(\SUMB[9][2] ), 
        .CO(\CARRYB[10][1] ), .S(\SUMB[10][1] ) );
  FADDX1 S2_10_2 ( .A(\ab[10][2] ), .B(\CARRYB[9][2] ), .CI(\SUMB[9][3] ), 
        .CO(\CARRYB[10][2] ), .S(\SUMB[10][2] ) );
  FADDX1 S2_10_3 ( .A(\ab[10][3] ), .B(\CARRYB[9][3] ), .CI(\SUMB[9][4] ), 
        .CO(\CARRYB[10][3] ), .S(\SUMB[10][3] ) );
  FADDX1 S2_10_4 ( .A(\ab[10][4] ), .B(\CARRYB[9][4] ), .CI(\SUMB[9][5] ), 
        .CO(\CARRYB[10][4] ), .S(\SUMB[10][4] ) );
  FADDX1 S2_10_5 ( .A(\ab[10][5] ), .B(\CARRYB[9][5] ), .CI(\SUMB[9][6] ), 
        .CO(\CARRYB[10][5] ), .S(\SUMB[10][5] ) );
  FADDX1 S2_10_6 ( .A(\ab[10][6] ), .B(\CARRYB[9][6] ), .CI(\SUMB[9][7] ), 
        .CO(\CARRYB[10][6] ), .S(\SUMB[10][6] ) );
  FADDX1 S2_10_7 ( .A(\ab[10][7] ), .B(\CARRYB[9][7] ), .CI(\SUMB[9][8] ), 
        .CO(\CARRYB[10][7] ), .S(\SUMB[10][7] ) );
  FADDX1 S2_10_8 ( .A(\ab[10][8] ), .B(\CARRYB[9][8] ), .CI(\SUMB[9][9] ), 
        .CO(\CARRYB[10][8] ), .S(\SUMB[10][8] ) );
  FADDX1 S2_10_9 ( .A(\ab[10][9] ), .B(\CARRYB[9][9] ), .CI(\SUMB[9][10] ), 
        .CO(\CARRYB[10][9] ), .S(\SUMB[10][9] ) );
  FADDX1 S2_10_10 ( .A(\ab[10][10] ), .B(\CARRYB[9][10] ), .CI(\SUMB[9][11] ), 
        .CO(\CARRYB[10][10] ), .S(\SUMB[10][10] ) );
  FADDX1 S2_10_11 ( .A(\ab[10][11] ), .B(\CARRYB[9][11] ), .CI(\SUMB[9][12] ), 
        .CO(\CARRYB[10][11] ), .S(\SUMB[10][11] ) );
  FADDX1 S2_10_12 ( .A(\ab[10][12] ), .B(\CARRYB[9][12] ), .CI(\SUMB[9][13] ), 
        .CO(\CARRYB[10][12] ), .S(\SUMB[10][12] ) );
  FADDX1 S2_10_13 ( .A(\ab[10][13] ), .B(\CARRYB[9][13] ), .CI(\SUMB[9][14] ), 
        .CO(\CARRYB[10][13] ), .S(\SUMB[10][13] ) );
  FADDX1 S2_10_14 ( .A(\ab[10][14] ), .B(\CARRYB[9][14] ), .CI(\SUMB[9][15] ), 
        .CO(\CARRYB[10][14] ), .S(\SUMB[10][14] ) );
  FADDX1 S2_10_15 ( .A(\ab[10][15] ), .B(\CARRYB[9][15] ), .CI(\SUMB[9][16] ), 
        .CO(\CARRYB[10][15] ), .S(\SUMB[10][15] ) );
  FADDX1 S2_10_16 ( .A(\ab[10][16] ), .B(\CARRYB[9][16] ), .CI(\SUMB[9][17] ), 
        .CO(\CARRYB[10][16] ), .S(\SUMB[10][16] ) );
  FADDX1 S2_10_17 ( .A(\ab[10][17] ), .B(\CARRYB[9][17] ), .CI(\SUMB[9][18] ), 
        .CO(\CARRYB[10][17] ), .S(\SUMB[10][17] ) );
  FADDX1 S2_10_18 ( .A(\ab[10][18] ), .B(\CARRYB[9][18] ), .CI(\SUMB[9][19] ), 
        .CO(\CARRYB[10][18] ), .S(\SUMB[10][18] ) );
  FADDX1 S2_10_19 ( .A(\ab[10][19] ), .B(\CARRYB[9][19] ), .CI(\SUMB[9][20] ), 
        .CO(\CARRYB[10][19] ), .S(\SUMB[10][19] ) );
  FADDX1 S2_10_20 ( .A(\ab[10][20] ), .B(\CARRYB[9][20] ), .CI(\SUMB[9][21] ), 
        .CO(\CARRYB[10][20] ), .S(\SUMB[10][20] ) );
  FADDX1 S2_10_21 ( .A(\ab[10][21] ), .B(\CARRYB[9][21] ), .CI(\SUMB[9][22] ), 
        .CO(\CARRYB[10][21] ), .S(\SUMB[10][21] ) );
  FADDX1 S3_10_22 ( .A(\ab[10][22] ), .B(\CARRYB[9][22] ), .CI(\ab[9][23] ), 
        .CO(\CARRYB[10][22] ), .S(\SUMB[10][22] ) );
  FADDX1 S1_9_0 ( .A(\ab[9][0] ), .B(\CARRYB[8][0] ), .CI(\SUMB[8][1] ), .CO(
        \CARRYB[9][0] ), .S(\A1[7] ) );
  FADDX1 S2_9_1 ( .A(\ab[9][1] ), .B(\CARRYB[8][1] ), .CI(\SUMB[8][2] ), .CO(
        \CARRYB[9][1] ), .S(\SUMB[9][1] ) );
  FADDX1 S2_9_2 ( .A(\ab[9][2] ), .B(\CARRYB[8][2] ), .CI(\SUMB[8][3] ), .CO(
        \CARRYB[9][2] ), .S(\SUMB[9][2] ) );
  FADDX1 S2_9_3 ( .A(\ab[9][3] ), .B(\CARRYB[8][3] ), .CI(\SUMB[8][4] ), .CO(
        \CARRYB[9][3] ), .S(\SUMB[9][3] ) );
  FADDX1 S2_9_4 ( .A(\ab[9][4] ), .B(\CARRYB[8][4] ), .CI(\SUMB[8][5] ), .CO(
        \CARRYB[9][4] ), .S(\SUMB[9][4] ) );
  FADDX1 S2_9_5 ( .A(\ab[9][5] ), .B(\CARRYB[8][5] ), .CI(\SUMB[8][6] ), .CO(
        \CARRYB[9][5] ), .S(\SUMB[9][5] ) );
  FADDX1 S2_9_6 ( .A(\ab[9][6] ), .B(\CARRYB[8][6] ), .CI(\SUMB[8][7] ), .CO(
        \CARRYB[9][6] ), .S(\SUMB[9][6] ) );
  FADDX1 S2_9_7 ( .A(\ab[9][7] ), .B(\CARRYB[8][7] ), .CI(\SUMB[8][8] ), .CO(
        \CARRYB[9][7] ), .S(\SUMB[9][7] ) );
  FADDX1 S2_9_8 ( .A(\ab[9][8] ), .B(\CARRYB[8][8] ), .CI(\SUMB[8][9] ), .CO(
        \CARRYB[9][8] ), .S(\SUMB[9][8] ) );
  FADDX1 S2_9_9 ( .A(\ab[9][9] ), .B(\CARRYB[8][9] ), .CI(\SUMB[8][10] ), .CO(
        \CARRYB[9][9] ), .S(\SUMB[9][9] ) );
  FADDX1 S2_9_10 ( .A(\ab[9][10] ), .B(\CARRYB[8][10] ), .CI(\SUMB[8][11] ), 
        .CO(\CARRYB[9][10] ), .S(\SUMB[9][10] ) );
  FADDX1 S2_9_11 ( .A(\ab[9][11] ), .B(\CARRYB[8][11] ), .CI(\SUMB[8][12] ), 
        .CO(\CARRYB[9][11] ), .S(\SUMB[9][11] ) );
  FADDX1 S2_9_12 ( .A(\ab[9][12] ), .B(\CARRYB[8][12] ), .CI(\SUMB[8][13] ), 
        .CO(\CARRYB[9][12] ), .S(\SUMB[9][12] ) );
  FADDX1 S2_9_13 ( .A(\ab[9][13] ), .B(\CARRYB[8][13] ), .CI(\SUMB[8][14] ), 
        .CO(\CARRYB[9][13] ), .S(\SUMB[9][13] ) );
  FADDX1 S2_9_14 ( .A(\ab[9][14] ), .B(\CARRYB[8][14] ), .CI(\SUMB[8][15] ), 
        .CO(\CARRYB[9][14] ), .S(\SUMB[9][14] ) );
  FADDX1 S2_9_15 ( .A(\ab[9][15] ), .B(\CARRYB[8][15] ), .CI(\SUMB[8][16] ), 
        .CO(\CARRYB[9][15] ), .S(\SUMB[9][15] ) );
  FADDX1 S2_9_16 ( .A(\ab[9][16] ), .B(\CARRYB[8][16] ), .CI(\SUMB[8][17] ), 
        .CO(\CARRYB[9][16] ), .S(\SUMB[9][16] ) );
  FADDX1 S2_9_17 ( .A(\ab[9][17] ), .B(\CARRYB[8][17] ), .CI(\SUMB[8][18] ), 
        .CO(\CARRYB[9][17] ), .S(\SUMB[9][17] ) );
  FADDX1 S2_9_18 ( .A(\ab[9][18] ), .B(\CARRYB[8][18] ), .CI(\SUMB[8][19] ), 
        .CO(\CARRYB[9][18] ), .S(\SUMB[9][18] ) );
  FADDX1 S2_9_19 ( .A(\ab[9][19] ), .B(\CARRYB[8][19] ), .CI(\SUMB[8][20] ), 
        .CO(\CARRYB[9][19] ), .S(\SUMB[9][19] ) );
  FADDX1 S2_9_20 ( .A(\ab[9][20] ), .B(\CARRYB[8][20] ), .CI(\SUMB[8][21] ), 
        .CO(\CARRYB[9][20] ), .S(\SUMB[9][20] ) );
  FADDX1 S2_9_21 ( .A(\ab[9][21] ), .B(\CARRYB[8][21] ), .CI(\SUMB[8][22] ), 
        .CO(\CARRYB[9][21] ), .S(\SUMB[9][21] ) );
  FADDX1 S3_9_22 ( .A(\ab[9][22] ), .B(\CARRYB[8][22] ), .CI(\ab[8][23] ), 
        .CO(\CARRYB[9][22] ), .S(\SUMB[9][22] ) );
  FADDX1 S1_8_0 ( .A(\ab[8][0] ), .B(\CARRYB[7][0] ), .CI(\SUMB[7][1] ), .CO(
        \CARRYB[8][0] ), .S(\A1[6] ) );
  FADDX1 S2_8_1 ( .A(\ab[8][1] ), .B(\CARRYB[7][1] ), .CI(\SUMB[7][2] ), .CO(
        \CARRYB[8][1] ), .S(\SUMB[8][1] ) );
  FADDX1 S2_8_2 ( .A(\ab[8][2] ), .B(\CARRYB[7][2] ), .CI(\SUMB[7][3] ), .CO(
        \CARRYB[8][2] ), .S(\SUMB[8][2] ) );
  FADDX1 S2_8_3 ( .A(\ab[8][3] ), .B(\CARRYB[7][3] ), .CI(\SUMB[7][4] ), .CO(
        \CARRYB[8][3] ), .S(\SUMB[8][3] ) );
  FADDX1 S2_8_4 ( .A(\ab[8][4] ), .B(\CARRYB[7][4] ), .CI(\SUMB[7][5] ), .CO(
        \CARRYB[8][4] ), .S(\SUMB[8][4] ) );
  FADDX1 S2_8_5 ( .A(\ab[8][5] ), .B(\CARRYB[7][5] ), .CI(\SUMB[7][6] ), .CO(
        \CARRYB[8][5] ), .S(\SUMB[8][5] ) );
  FADDX1 S2_8_6 ( .A(\ab[8][6] ), .B(\CARRYB[7][6] ), .CI(\SUMB[7][7] ), .CO(
        \CARRYB[8][6] ), .S(\SUMB[8][6] ) );
  FADDX1 S2_8_7 ( .A(\ab[8][7] ), .B(\CARRYB[7][7] ), .CI(\SUMB[7][8] ), .CO(
        \CARRYB[8][7] ), .S(\SUMB[8][7] ) );
  FADDX1 S2_8_8 ( .A(\ab[8][8] ), .B(\CARRYB[7][8] ), .CI(\SUMB[7][9] ), .CO(
        \CARRYB[8][8] ), .S(\SUMB[8][8] ) );
  FADDX1 S2_8_9 ( .A(\ab[8][9] ), .B(\CARRYB[7][9] ), .CI(\SUMB[7][10] ), .CO(
        \CARRYB[8][9] ), .S(\SUMB[8][9] ) );
  FADDX1 S2_8_10 ( .A(\ab[8][10] ), .B(\CARRYB[7][10] ), .CI(\SUMB[7][11] ), 
        .CO(\CARRYB[8][10] ), .S(\SUMB[8][10] ) );
  FADDX1 S2_8_11 ( .A(\ab[8][11] ), .B(\CARRYB[7][11] ), .CI(\SUMB[7][12] ), 
        .CO(\CARRYB[8][11] ), .S(\SUMB[8][11] ) );
  FADDX1 S2_8_12 ( .A(\ab[8][12] ), .B(\CARRYB[7][12] ), .CI(\SUMB[7][13] ), 
        .CO(\CARRYB[8][12] ), .S(\SUMB[8][12] ) );
  FADDX1 S2_8_13 ( .A(\ab[8][13] ), .B(\CARRYB[7][13] ), .CI(\SUMB[7][14] ), 
        .CO(\CARRYB[8][13] ), .S(\SUMB[8][13] ) );
  FADDX1 S2_8_14 ( .A(\ab[8][14] ), .B(\CARRYB[7][14] ), .CI(\SUMB[7][15] ), 
        .CO(\CARRYB[8][14] ), .S(\SUMB[8][14] ) );
  FADDX1 S2_8_15 ( .A(\ab[8][15] ), .B(\CARRYB[7][15] ), .CI(\SUMB[7][16] ), 
        .CO(\CARRYB[8][15] ), .S(\SUMB[8][15] ) );
  FADDX1 S2_8_16 ( .A(\ab[8][16] ), .B(\CARRYB[7][16] ), .CI(\SUMB[7][17] ), 
        .CO(\CARRYB[8][16] ), .S(\SUMB[8][16] ) );
  FADDX1 S2_8_17 ( .A(\ab[8][17] ), .B(\CARRYB[7][17] ), .CI(\SUMB[7][18] ), 
        .CO(\CARRYB[8][17] ), .S(\SUMB[8][17] ) );
  FADDX1 S2_8_18 ( .A(\ab[8][18] ), .B(\CARRYB[7][18] ), .CI(\SUMB[7][19] ), 
        .CO(\CARRYB[8][18] ), .S(\SUMB[8][18] ) );
  FADDX1 S2_8_19 ( .A(\ab[8][19] ), .B(\CARRYB[7][19] ), .CI(\SUMB[7][20] ), 
        .CO(\CARRYB[8][19] ), .S(\SUMB[8][19] ) );
  FADDX1 S2_8_20 ( .A(\ab[8][20] ), .B(\CARRYB[7][20] ), .CI(\SUMB[7][21] ), 
        .CO(\CARRYB[8][20] ), .S(\SUMB[8][20] ) );
  FADDX1 S2_8_21 ( .A(\ab[8][21] ), .B(\CARRYB[7][21] ), .CI(\SUMB[7][22] ), 
        .CO(\CARRYB[8][21] ), .S(\SUMB[8][21] ) );
  FADDX1 S3_8_22 ( .A(\ab[8][22] ), .B(\CARRYB[7][22] ), .CI(\ab[7][23] ), 
        .CO(\CARRYB[8][22] ), .S(\SUMB[8][22] ) );
  FADDX1 S1_7_0 ( .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .CI(\SUMB[6][1] ), .CO(
        \CARRYB[7][0] ), .S(\A1[5] ) );
  FADDX1 S2_7_1 ( .A(\ab[7][1] ), .B(\CARRYB[6][1] ), .CI(\SUMB[6][2] ), .CO(
        \CARRYB[7][1] ), .S(\SUMB[7][1] ) );
  FADDX1 S2_7_2 ( .A(\ab[7][2] ), .B(\CARRYB[6][2] ), .CI(\SUMB[6][3] ), .CO(
        \CARRYB[7][2] ), .S(\SUMB[7][2] ) );
  FADDX1 S2_7_3 ( .A(\ab[7][3] ), .B(\CARRYB[6][3] ), .CI(\SUMB[6][4] ), .CO(
        \CARRYB[7][3] ), .S(\SUMB[7][3] ) );
  FADDX1 S2_7_4 ( .A(\ab[7][4] ), .B(\CARRYB[6][4] ), .CI(\SUMB[6][5] ), .CO(
        \CARRYB[7][4] ), .S(\SUMB[7][4] ) );
  FADDX1 S2_7_5 ( .A(\ab[7][5] ), .B(\CARRYB[6][5] ), .CI(\SUMB[6][6] ), .CO(
        \CARRYB[7][5] ), .S(\SUMB[7][5] ) );
  FADDX1 S2_7_6 ( .A(\ab[7][6] ), .B(\CARRYB[6][6] ), .CI(\SUMB[6][7] ), .CO(
        \CARRYB[7][6] ), .S(\SUMB[7][6] ) );
  FADDX1 S2_7_7 ( .A(\ab[7][7] ), .B(\CARRYB[6][7] ), .CI(\SUMB[6][8] ), .CO(
        \CARRYB[7][7] ), .S(\SUMB[7][7] ) );
  FADDX1 S2_7_8 ( .A(\ab[7][8] ), .B(\CARRYB[6][8] ), .CI(\SUMB[6][9] ), .CO(
        \CARRYB[7][8] ), .S(\SUMB[7][8] ) );
  FADDX1 S2_7_9 ( .A(\ab[7][9] ), .B(\CARRYB[6][9] ), .CI(\SUMB[6][10] ), .CO(
        \CARRYB[7][9] ), .S(\SUMB[7][9] ) );
  FADDX1 S2_7_10 ( .A(\ab[7][10] ), .B(\CARRYB[6][10] ), .CI(\SUMB[6][11] ), 
        .CO(\CARRYB[7][10] ), .S(\SUMB[7][10] ) );
  FADDX1 S2_7_11 ( .A(\ab[7][11] ), .B(\CARRYB[6][11] ), .CI(\SUMB[6][12] ), 
        .CO(\CARRYB[7][11] ), .S(\SUMB[7][11] ) );
  FADDX1 S2_7_12 ( .A(\ab[7][12] ), .B(\CARRYB[6][12] ), .CI(\SUMB[6][13] ), 
        .CO(\CARRYB[7][12] ), .S(\SUMB[7][12] ) );
  FADDX1 S2_7_13 ( .A(\ab[7][13] ), .B(\CARRYB[6][13] ), .CI(\SUMB[6][14] ), 
        .CO(\CARRYB[7][13] ), .S(\SUMB[7][13] ) );
  FADDX1 S2_7_14 ( .A(\ab[7][14] ), .B(\CARRYB[6][14] ), .CI(\SUMB[6][15] ), 
        .CO(\CARRYB[7][14] ), .S(\SUMB[7][14] ) );
  FADDX1 S2_7_15 ( .A(\ab[7][15] ), .B(\CARRYB[6][15] ), .CI(\SUMB[6][16] ), 
        .CO(\CARRYB[7][15] ), .S(\SUMB[7][15] ) );
  FADDX1 S2_7_16 ( .A(\ab[7][16] ), .B(\CARRYB[6][16] ), .CI(\SUMB[6][17] ), 
        .CO(\CARRYB[7][16] ), .S(\SUMB[7][16] ) );
  FADDX1 S2_7_17 ( .A(\ab[7][17] ), .B(\CARRYB[6][17] ), .CI(\SUMB[6][18] ), 
        .CO(\CARRYB[7][17] ), .S(\SUMB[7][17] ) );
  FADDX1 S2_7_18 ( .A(\ab[7][18] ), .B(\CARRYB[6][18] ), .CI(\SUMB[6][19] ), 
        .CO(\CARRYB[7][18] ), .S(\SUMB[7][18] ) );
  FADDX1 S2_7_19 ( .A(\ab[7][19] ), .B(\CARRYB[6][19] ), .CI(\SUMB[6][20] ), 
        .CO(\CARRYB[7][19] ), .S(\SUMB[7][19] ) );
  FADDX1 S2_7_20 ( .A(\ab[7][20] ), .B(\CARRYB[6][20] ), .CI(\SUMB[6][21] ), 
        .CO(\CARRYB[7][20] ), .S(\SUMB[7][20] ) );
  FADDX1 S2_7_21 ( .A(\ab[7][21] ), .B(\CARRYB[6][21] ), .CI(\SUMB[6][22] ), 
        .CO(\CARRYB[7][21] ), .S(\SUMB[7][21] ) );
  FADDX1 S3_7_22 ( .A(\ab[7][22] ), .B(\CARRYB[6][22] ), .CI(\ab[6][23] ), 
        .CO(\CARRYB[7][22] ), .S(\SUMB[7][22] ) );
  FADDX1 S1_6_0 ( .A(\ab[6][0] ), .B(\CARRYB[5][0] ), .CI(\SUMB[5][1] ), .CO(
        \CARRYB[6][0] ), .S(\A1[4] ) );
  FADDX1 S2_6_1 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .CI(\SUMB[5][2] ), .CO(
        \CARRYB[6][1] ), .S(\SUMB[6][1] ) );
  FADDX1 S2_6_2 ( .A(\ab[6][2] ), .B(\CARRYB[5][2] ), .CI(\SUMB[5][3] ), .CO(
        \CARRYB[6][2] ), .S(\SUMB[6][2] ) );
  FADDX1 S2_6_3 ( .A(\ab[6][3] ), .B(\CARRYB[5][3] ), .CI(\SUMB[5][4] ), .CO(
        \CARRYB[6][3] ), .S(\SUMB[6][3] ) );
  FADDX1 S2_6_4 ( .A(\ab[6][4] ), .B(\CARRYB[5][4] ), .CI(\SUMB[5][5] ), .CO(
        \CARRYB[6][4] ), .S(\SUMB[6][4] ) );
  FADDX1 S2_6_5 ( .A(\ab[6][5] ), .B(\CARRYB[5][5] ), .CI(\SUMB[5][6] ), .CO(
        \CARRYB[6][5] ), .S(\SUMB[6][5] ) );
  FADDX1 S2_6_6 ( .A(\ab[6][6] ), .B(\CARRYB[5][6] ), .CI(\SUMB[5][7] ), .CO(
        \CARRYB[6][6] ), .S(\SUMB[6][6] ) );
  FADDX1 S2_6_7 ( .A(\ab[6][7] ), .B(\CARRYB[5][7] ), .CI(\SUMB[5][8] ), .CO(
        \CARRYB[6][7] ), .S(\SUMB[6][7] ) );
  FADDX1 S2_6_8 ( .A(\ab[6][8] ), .B(\CARRYB[5][8] ), .CI(\SUMB[5][9] ), .CO(
        \CARRYB[6][8] ), .S(\SUMB[6][8] ) );
  FADDX1 S2_6_9 ( .A(\ab[6][9] ), .B(\CARRYB[5][9] ), .CI(\SUMB[5][10] ), .CO(
        \CARRYB[6][9] ), .S(\SUMB[6][9] ) );
  FADDX1 S2_6_10 ( .A(\ab[6][10] ), .B(\CARRYB[5][10] ), .CI(\SUMB[5][11] ), 
        .CO(\CARRYB[6][10] ), .S(\SUMB[6][10] ) );
  FADDX1 S2_6_11 ( .A(\ab[6][11] ), .B(\CARRYB[5][11] ), .CI(\SUMB[5][12] ), 
        .CO(\CARRYB[6][11] ), .S(\SUMB[6][11] ) );
  FADDX1 S2_6_12 ( .A(\ab[6][12] ), .B(\CARRYB[5][12] ), .CI(\SUMB[5][13] ), 
        .CO(\CARRYB[6][12] ), .S(\SUMB[6][12] ) );
  FADDX1 S2_6_13 ( .A(\ab[6][13] ), .B(\CARRYB[5][13] ), .CI(\SUMB[5][14] ), 
        .CO(\CARRYB[6][13] ), .S(\SUMB[6][13] ) );
  FADDX1 S2_6_14 ( .A(\ab[6][14] ), .B(\CARRYB[5][14] ), .CI(\SUMB[5][15] ), 
        .CO(\CARRYB[6][14] ), .S(\SUMB[6][14] ) );
  FADDX1 S2_6_15 ( .A(\ab[6][15] ), .B(\CARRYB[5][15] ), .CI(\SUMB[5][16] ), 
        .CO(\CARRYB[6][15] ), .S(\SUMB[6][15] ) );
  FADDX1 S2_6_16 ( .A(\ab[6][16] ), .B(\CARRYB[5][16] ), .CI(\SUMB[5][17] ), 
        .CO(\CARRYB[6][16] ), .S(\SUMB[6][16] ) );
  FADDX1 S2_6_17 ( .A(\ab[6][17] ), .B(\CARRYB[5][17] ), .CI(\SUMB[5][18] ), 
        .CO(\CARRYB[6][17] ), .S(\SUMB[6][17] ) );
  FADDX1 S2_6_18 ( .A(\ab[6][18] ), .B(\CARRYB[5][18] ), .CI(\SUMB[5][19] ), 
        .CO(\CARRYB[6][18] ), .S(\SUMB[6][18] ) );
  FADDX1 S2_6_19 ( .A(\ab[6][19] ), .B(\CARRYB[5][19] ), .CI(\SUMB[5][20] ), 
        .CO(\CARRYB[6][19] ), .S(\SUMB[6][19] ) );
  FADDX1 S2_6_20 ( .A(\ab[6][20] ), .B(\CARRYB[5][20] ), .CI(\SUMB[5][21] ), 
        .CO(\CARRYB[6][20] ), .S(\SUMB[6][20] ) );
  FADDX1 S2_6_21 ( .A(\ab[6][21] ), .B(\CARRYB[5][21] ), .CI(\SUMB[5][22] ), 
        .CO(\CARRYB[6][21] ), .S(\SUMB[6][21] ) );
  FADDX1 S3_6_22 ( .A(\ab[6][22] ), .B(\CARRYB[5][22] ), .CI(\ab[5][23] ), 
        .CO(\CARRYB[6][22] ), .S(\SUMB[6][22] ) );
  FADDX1 S1_5_0 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .CI(\SUMB[4][1] ), .CO(
        \CARRYB[5][0] ), .S(\A1[3] ) );
  FADDX1 S2_5_1 ( .A(\ab[5][1] ), .B(\CARRYB[4][1] ), .CI(\SUMB[4][2] ), .CO(
        \CARRYB[5][1] ), .S(\SUMB[5][1] ) );
  FADDX1 S2_5_2 ( .A(\ab[5][2] ), .B(\CARRYB[4][2] ), .CI(\SUMB[4][3] ), .CO(
        \CARRYB[5][2] ), .S(\SUMB[5][2] ) );
  FADDX1 S2_5_3 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .CI(\SUMB[4][4] ), .CO(
        \CARRYB[5][3] ), .S(\SUMB[5][3] ) );
  FADDX1 S2_5_4 ( .A(\ab[5][4] ), .B(\CARRYB[4][4] ), .CI(\SUMB[4][5] ), .CO(
        \CARRYB[5][4] ), .S(\SUMB[5][4] ) );
  FADDX1 S2_5_5 ( .A(\ab[5][5] ), .B(\CARRYB[4][5] ), .CI(\SUMB[4][6] ), .CO(
        \CARRYB[5][5] ), .S(\SUMB[5][5] ) );
  FADDX1 S2_5_6 ( .A(\ab[5][6] ), .B(\CARRYB[4][6] ), .CI(\SUMB[4][7] ), .CO(
        \CARRYB[5][6] ), .S(\SUMB[5][6] ) );
  FADDX1 S2_5_7 ( .A(\ab[5][7] ), .B(\CARRYB[4][7] ), .CI(\SUMB[4][8] ), .CO(
        \CARRYB[5][7] ), .S(\SUMB[5][7] ) );
  FADDX1 S2_5_8 ( .A(\ab[5][8] ), .B(\CARRYB[4][8] ), .CI(\SUMB[4][9] ), .CO(
        \CARRYB[5][8] ), .S(\SUMB[5][8] ) );
  FADDX1 S2_5_9 ( .A(\ab[5][9] ), .B(\CARRYB[4][9] ), .CI(\SUMB[4][10] ), .CO(
        \CARRYB[5][9] ), .S(\SUMB[5][9] ) );
  FADDX1 S2_5_10 ( .A(\ab[5][10] ), .B(\CARRYB[4][10] ), .CI(\SUMB[4][11] ), 
        .CO(\CARRYB[5][10] ), .S(\SUMB[5][10] ) );
  FADDX1 S2_5_11 ( .A(\ab[5][11] ), .B(\CARRYB[4][11] ), .CI(\SUMB[4][12] ), 
        .CO(\CARRYB[5][11] ), .S(\SUMB[5][11] ) );
  FADDX1 S2_5_12 ( .A(\ab[5][12] ), .B(\CARRYB[4][12] ), .CI(\SUMB[4][13] ), 
        .CO(\CARRYB[5][12] ), .S(\SUMB[5][12] ) );
  FADDX1 S2_5_13 ( .A(\ab[5][13] ), .B(\CARRYB[4][13] ), .CI(\SUMB[4][14] ), 
        .CO(\CARRYB[5][13] ), .S(\SUMB[5][13] ) );
  FADDX1 S2_5_14 ( .A(\ab[5][14] ), .B(\CARRYB[4][14] ), .CI(\SUMB[4][15] ), 
        .CO(\CARRYB[5][14] ), .S(\SUMB[5][14] ) );
  FADDX1 S2_5_15 ( .A(\ab[5][15] ), .B(\CARRYB[4][15] ), .CI(\SUMB[4][16] ), 
        .CO(\CARRYB[5][15] ), .S(\SUMB[5][15] ) );
  FADDX1 S2_5_16 ( .A(\ab[5][16] ), .B(\CARRYB[4][16] ), .CI(\SUMB[4][17] ), 
        .CO(\CARRYB[5][16] ), .S(\SUMB[5][16] ) );
  FADDX1 S2_5_17 ( .A(\ab[5][17] ), .B(\CARRYB[4][17] ), .CI(\SUMB[4][18] ), 
        .CO(\CARRYB[5][17] ), .S(\SUMB[5][17] ) );
  FADDX1 S2_5_18 ( .A(\ab[5][18] ), .B(\CARRYB[4][18] ), .CI(\SUMB[4][19] ), 
        .CO(\CARRYB[5][18] ), .S(\SUMB[5][18] ) );
  FADDX1 S2_5_19 ( .A(\ab[5][19] ), .B(\CARRYB[4][19] ), .CI(\SUMB[4][20] ), 
        .CO(\CARRYB[5][19] ), .S(\SUMB[5][19] ) );
  FADDX1 S2_5_20 ( .A(\ab[5][20] ), .B(\CARRYB[4][20] ), .CI(\SUMB[4][21] ), 
        .CO(\CARRYB[5][20] ), .S(\SUMB[5][20] ) );
  FADDX1 S2_5_21 ( .A(\ab[5][21] ), .B(\CARRYB[4][21] ), .CI(\SUMB[4][22] ), 
        .CO(\CARRYB[5][21] ), .S(\SUMB[5][21] ) );
  FADDX1 S3_5_22 ( .A(\ab[5][22] ), .B(\CARRYB[4][22] ), .CI(\ab[4][23] ), 
        .CO(\CARRYB[5][22] ), .S(\SUMB[5][22] ) );
  FADDX1 S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .CI(\SUMB[3][1] ), .CO(
        \CARRYB[4][0] ), .S(\A1[2] ) );
  FADDX1 S2_4_1 ( .A(\ab[4][1] ), .B(\CARRYB[3][1] ), .CI(\SUMB[3][2] ), .CO(
        \CARRYB[4][1] ), .S(\SUMB[4][1] ) );
  FADDX1 S2_4_2 ( .A(\ab[4][2] ), .B(\CARRYB[3][2] ), .CI(\SUMB[3][3] ), .CO(
        \CARRYB[4][2] ), .S(\SUMB[4][2] ) );
  FADDX1 S2_4_3 ( .A(\ab[4][3] ), .B(\CARRYB[3][3] ), .CI(\SUMB[3][4] ), .CO(
        \CARRYB[4][3] ), .S(\SUMB[4][3] ) );
  FADDX1 S2_4_4 ( .A(\ab[4][4] ), .B(\CARRYB[3][4] ), .CI(\SUMB[3][5] ), .CO(
        \CARRYB[4][4] ), .S(\SUMB[4][4] ) );
  FADDX1 S2_4_5 ( .A(\ab[4][5] ), .B(\CARRYB[3][5] ), .CI(\SUMB[3][6] ), .CO(
        \CARRYB[4][5] ), .S(\SUMB[4][5] ) );
  FADDX1 S2_4_6 ( .A(\ab[4][6] ), .B(\CARRYB[3][6] ), .CI(\SUMB[3][7] ), .CO(
        \CARRYB[4][6] ), .S(\SUMB[4][6] ) );
  FADDX1 S2_4_7 ( .A(\ab[4][7] ), .B(\CARRYB[3][7] ), .CI(\SUMB[3][8] ), .CO(
        \CARRYB[4][7] ), .S(\SUMB[4][7] ) );
  FADDX1 S2_4_8 ( .A(\ab[4][8] ), .B(\CARRYB[3][8] ), .CI(\SUMB[3][9] ), .CO(
        \CARRYB[4][8] ), .S(\SUMB[4][8] ) );
  FADDX1 S2_4_9 ( .A(\ab[4][9] ), .B(\CARRYB[3][9] ), .CI(\SUMB[3][10] ), .CO(
        \CARRYB[4][9] ), .S(\SUMB[4][9] ) );
  FADDX1 S2_4_10 ( .A(\ab[4][10] ), .B(\CARRYB[3][10] ), .CI(\SUMB[3][11] ), 
        .CO(\CARRYB[4][10] ), .S(\SUMB[4][10] ) );
  FADDX1 S2_4_11 ( .A(\ab[4][11] ), .B(\CARRYB[3][11] ), .CI(\SUMB[3][12] ), 
        .CO(\CARRYB[4][11] ), .S(\SUMB[4][11] ) );
  FADDX1 S2_4_12 ( .A(\ab[4][12] ), .B(\CARRYB[3][12] ), .CI(\SUMB[3][13] ), 
        .CO(\CARRYB[4][12] ), .S(\SUMB[4][12] ) );
  FADDX1 S2_4_13 ( .A(\ab[4][13] ), .B(\CARRYB[3][13] ), .CI(\SUMB[3][14] ), 
        .CO(\CARRYB[4][13] ), .S(\SUMB[4][13] ) );
  FADDX1 S2_4_14 ( .A(\ab[4][14] ), .B(\CARRYB[3][14] ), .CI(\SUMB[3][15] ), 
        .CO(\CARRYB[4][14] ), .S(\SUMB[4][14] ) );
  FADDX1 S2_4_15 ( .A(\ab[4][15] ), .B(\CARRYB[3][15] ), .CI(\SUMB[3][16] ), 
        .CO(\CARRYB[4][15] ), .S(\SUMB[4][15] ) );
  FADDX1 S2_4_16 ( .A(\ab[4][16] ), .B(\CARRYB[3][16] ), .CI(\SUMB[3][17] ), 
        .CO(\CARRYB[4][16] ), .S(\SUMB[4][16] ) );
  FADDX1 S2_4_17 ( .A(\ab[4][17] ), .B(\CARRYB[3][17] ), .CI(\SUMB[3][18] ), 
        .CO(\CARRYB[4][17] ), .S(\SUMB[4][17] ) );
  FADDX1 S2_4_18 ( .A(\ab[4][18] ), .B(\CARRYB[3][18] ), .CI(\SUMB[3][19] ), 
        .CO(\CARRYB[4][18] ), .S(\SUMB[4][18] ) );
  FADDX1 S2_4_19 ( .A(\ab[4][19] ), .B(\CARRYB[3][19] ), .CI(\SUMB[3][20] ), 
        .CO(\CARRYB[4][19] ), .S(\SUMB[4][19] ) );
  FADDX1 S2_4_20 ( .A(\ab[4][20] ), .B(\CARRYB[3][20] ), .CI(\SUMB[3][21] ), 
        .CO(\CARRYB[4][20] ), .S(\SUMB[4][20] ) );
  FADDX1 S2_4_21 ( .A(\ab[4][21] ), .B(\CARRYB[3][21] ), .CI(\SUMB[3][22] ), 
        .CO(\CARRYB[4][21] ), .S(\SUMB[4][21] ) );
  FADDX1 S3_4_22 ( .A(\ab[4][22] ), .B(\CARRYB[3][22] ), .CI(\ab[3][23] ), 
        .CO(\CARRYB[4][22] ), .S(\SUMB[4][22] ) );
  FADDX1 S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .CI(\SUMB[2][1] ), .CO(
        \CARRYB[3][0] ), .S(\A1[1] ) );
  FADDX1 S2_3_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .CI(\SUMB[2][2] ), .CO(
        \CARRYB[3][1] ), .S(\SUMB[3][1] ) );
  FADDX1 S2_3_2 ( .A(\ab[3][2] ), .B(\CARRYB[2][2] ), .CI(\SUMB[2][3] ), .CO(
        \CARRYB[3][2] ), .S(\SUMB[3][2] ) );
  FADDX1 S2_3_3 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .CI(\SUMB[2][4] ), .CO(
        \CARRYB[3][3] ), .S(\SUMB[3][3] ) );
  FADDX1 S2_3_4 ( .A(\ab[3][4] ), .B(\CARRYB[2][4] ), .CI(\SUMB[2][5] ), .CO(
        \CARRYB[3][4] ), .S(\SUMB[3][4] ) );
  FADDX1 S2_3_5 ( .A(\ab[3][5] ), .B(\CARRYB[2][5] ), .CI(\SUMB[2][6] ), .CO(
        \CARRYB[3][5] ), .S(\SUMB[3][5] ) );
  FADDX1 S2_3_6 ( .A(\ab[3][6] ), .B(\CARRYB[2][6] ), .CI(\SUMB[2][7] ), .CO(
        \CARRYB[3][6] ), .S(\SUMB[3][6] ) );
  FADDX1 S2_3_7 ( .A(\ab[3][7] ), .B(\CARRYB[2][7] ), .CI(\SUMB[2][8] ), .CO(
        \CARRYB[3][7] ), .S(\SUMB[3][7] ) );
  FADDX1 S2_3_8 ( .A(\ab[3][8] ), .B(\CARRYB[2][8] ), .CI(\SUMB[2][9] ), .CO(
        \CARRYB[3][8] ), .S(\SUMB[3][8] ) );
  FADDX1 S2_3_9 ( .A(\ab[3][9] ), .B(\CARRYB[2][9] ), .CI(\SUMB[2][10] ), .CO(
        \CARRYB[3][9] ), .S(\SUMB[3][9] ) );
  FADDX1 S2_3_10 ( .A(\ab[3][10] ), .B(\CARRYB[2][10] ), .CI(\SUMB[2][11] ), 
        .CO(\CARRYB[3][10] ), .S(\SUMB[3][10] ) );
  FADDX1 S2_3_11 ( .A(\ab[3][11] ), .B(\CARRYB[2][11] ), .CI(\SUMB[2][12] ), 
        .CO(\CARRYB[3][11] ), .S(\SUMB[3][11] ) );
  FADDX1 S2_3_12 ( .A(\ab[3][12] ), .B(\CARRYB[2][12] ), .CI(\SUMB[2][13] ), 
        .CO(\CARRYB[3][12] ), .S(\SUMB[3][12] ) );
  FADDX1 S2_3_13 ( .A(\ab[3][13] ), .B(\CARRYB[2][13] ), .CI(\SUMB[2][14] ), 
        .CO(\CARRYB[3][13] ), .S(\SUMB[3][13] ) );
  FADDX1 S2_3_14 ( .A(\ab[3][14] ), .B(\CARRYB[2][14] ), .CI(\SUMB[2][15] ), 
        .CO(\CARRYB[3][14] ), .S(\SUMB[3][14] ) );
  FADDX1 S2_3_15 ( .A(\ab[3][15] ), .B(\CARRYB[2][15] ), .CI(\SUMB[2][16] ), 
        .CO(\CARRYB[3][15] ), .S(\SUMB[3][15] ) );
  FADDX1 S2_3_16 ( .A(\ab[3][16] ), .B(\CARRYB[2][16] ), .CI(\SUMB[2][17] ), 
        .CO(\CARRYB[3][16] ), .S(\SUMB[3][16] ) );
  FADDX1 S2_3_17 ( .A(\ab[3][17] ), .B(\CARRYB[2][17] ), .CI(\SUMB[2][18] ), 
        .CO(\CARRYB[3][17] ), .S(\SUMB[3][17] ) );
  FADDX1 S2_3_18 ( .A(\ab[3][18] ), .B(\CARRYB[2][18] ), .CI(\SUMB[2][19] ), 
        .CO(\CARRYB[3][18] ), .S(\SUMB[3][18] ) );
  FADDX1 S2_3_19 ( .A(\ab[3][19] ), .B(\CARRYB[2][19] ), .CI(\SUMB[2][20] ), 
        .CO(\CARRYB[3][19] ), .S(\SUMB[3][19] ) );
  FADDX1 S2_3_20 ( .A(\ab[3][20] ), .B(\CARRYB[2][20] ), .CI(\SUMB[2][21] ), 
        .CO(\CARRYB[3][20] ), .S(\SUMB[3][20] ) );
  FADDX1 S2_3_21 ( .A(\ab[3][21] ), .B(\CARRYB[2][21] ), .CI(\SUMB[2][22] ), 
        .CO(\CARRYB[3][21] ), .S(\SUMB[3][21] ) );
  FADDX1 S3_3_22 ( .A(\ab[3][22] ), .B(\CARRYB[2][22] ), .CI(\ab[2][23] ), 
        .CO(\CARRYB[3][22] ), .S(\SUMB[3][22] ) );
  FADDX1 S1_2_0 ( .A(\ab[2][0] ), .B(\CARRYB[1][0] ), .CI(\SUMB[1][1] ), .CO(
        \CARRYB[2][0] ), .S(\A1[0] ) );
  FADDX1 S2_2_1 ( .A(\ab[2][1] ), .B(n3), .CI(\SUMB[1][2] ), .CO(
        \CARRYB[2][1] ), .S(\SUMB[2][1] ) );
  FADDX1 S2_2_2 ( .A(\ab[2][2] ), .B(n24), .CI(\SUMB[1][3] ), .CO(
        \CARRYB[2][2] ), .S(\SUMB[2][2] ) );
  FADDX1 S2_2_3 ( .A(\ab[2][3] ), .B(n23), .CI(\SUMB[1][4] ), .CO(
        \CARRYB[2][3] ), .S(\SUMB[2][3] ) );
  FADDX1 S2_2_4 ( .A(\ab[2][4] ), .B(n22), .CI(\SUMB[1][5] ), .CO(
        \CARRYB[2][4] ), .S(\SUMB[2][4] ) );
  FADDX1 S2_2_5 ( .A(\ab[2][5] ), .B(n21), .CI(\SUMB[1][6] ), .CO(
        \CARRYB[2][5] ), .S(\SUMB[2][5] ) );
  FADDX1 S2_2_6 ( .A(\ab[2][6] ), .B(n20), .CI(\SUMB[1][7] ), .CO(
        \CARRYB[2][6] ), .S(\SUMB[2][6] ) );
  FADDX1 S2_2_7 ( .A(\ab[2][7] ), .B(n19), .CI(\SUMB[1][8] ), .CO(
        \CARRYB[2][7] ), .S(\SUMB[2][7] ) );
  FADDX1 S2_2_8 ( .A(\ab[2][8] ), .B(n18), .CI(\SUMB[1][9] ), .CO(
        \CARRYB[2][8] ), .S(\SUMB[2][8] ) );
  FADDX1 S2_2_9 ( .A(\ab[2][9] ), .B(n17), .CI(\SUMB[1][10] ), .CO(
        \CARRYB[2][9] ), .S(\SUMB[2][9] ) );
  FADDX1 S2_2_10 ( .A(\ab[2][10] ), .B(n16), .CI(\SUMB[1][11] ), .CO(
        \CARRYB[2][10] ), .S(\SUMB[2][10] ) );
  FADDX1 S2_2_11 ( .A(\ab[2][11] ), .B(n15), .CI(\SUMB[1][12] ), .CO(
        \CARRYB[2][11] ), .S(\SUMB[2][11] ) );
  FADDX1 S2_2_12 ( .A(\ab[2][12] ), .B(n14), .CI(\SUMB[1][13] ), .CO(
        \CARRYB[2][12] ), .S(\SUMB[2][12] ) );
  FADDX1 S2_2_13 ( .A(\ab[2][13] ), .B(n13), .CI(\SUMB[1][14] ), .CO(
        \CARRYB[2][13] ), .S(\SUMB[2][13] ) );
  FADDX1 S2_2_14 ( .A(\ab[2][14] ), .B(n12), .CI(\SUMB[1][15] ), .CO(
        \CARRYB[2][14] ), .S(\SUMB[2][14] ) );
  FADDX1 S2_2_15 ( .A(\ab[2][15] ), .B(n11), .CI(\SUMB[1][16] ), .CO(
        \CARRYB[2][15] ), .S(\SUMB[2][15] ) );
  FADDX1 S2_2_16 ( .A(\ab[2][16] ), .B(n10), .CI(\SUMB[1][17] ), .CO(
        \CARRYB[2][16] ), .S(\SUMB[2][16] ) );
  FADDX1 S2_2_17 ( .A(\ab[2][17] ), .B(n9), .CI(\SUMB[1][18] ), .CO(
        \CARRYB[2][17] ), .S(\SUMB[2][17] ) );
  FADDX1 S2_2_18 ( .A(\ab[2][18] ), .B(n8), .CI(\SUMB[1][19] ), .CO(
        \CARRYB[2][18] ), .S(\SUMB[2][18] ) );
  FADDX1 S2_2_19 ( .A(\ab[2][19] ), .B(n7), .CI(\SUMB[1][20] ), .CO(
        \CARRYB[2][19] ), .S(\SUMB[2][19] ) );
  FADDX1 S2_2_20 ( .A(\ab[2][20] ), .B(n6), .CI(\SUMB[1][21] ), .CO(
        \CARRYB[2][20] ), .S(\SUMB[2][20] ) );
  FADDX1 S2_2_21 ( .A(\ab[2][21] ), .B(n5), .CI(\SUMB[1][22] ), .CO(
        \CARRYB[2][21] ), .S(\SUMB[2][21] ) );
  FADDX1 S3_2_22 ( .A(\ab[2][22] ), .B(n4), .CI(\ab[1][23] ), .CO(
        \CARRYB[2][22] ), .S(\SUMB[2][22] ) );
  fpalu_multiplier_DW01_add_1 FS_1 ( .A({1'b0, \A1[44] , \A1[43] , \A1[42] , 
        \A1[41] , \A1[40] , \A1[39] , \A1[38] , \A1[37] , \A1[36] , \A1[35] , 
        \A1[34] , \A1[33] , \A1[32] , \A1[31] , \A1[30] , \A1[29] , \A1[28] , 
        \A1[27] , \A1[26] , \A1[25] , \A1[24] , \A1[23] , \A1[22] , 
        \SUMB[23][0] , \A1[20] , \A1[19] , \A1[18] , \A1[17] , \A1[16] , 
        \A1[15] , \A1[14] , \A1[13] , \A1[12] , \A1[11] , \A1[10] , \A1[9] , 
        \A1[8] , \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] , 
        \A1[0] }), .B({n25, n26, n37, n36, n35, n34, n33, n32, n31, n30, n29, 
        n28, n27, n45, n44, n43, n42, n41, n40, n39, n38, n46, n47, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), 
        .SUM({PRODUCT[47:23], SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20}) );
  AND2X1 U2 ( .IN1(\ab[1][1] ), .IN2(\ab[0][2] ), .Q(n3) );
  AND2X1 U3 ( .IN1(\ab[1][22] ), .IN2(\ab[0][23] ), .Q(n4) );
  AND2X1 U4 ( .IN1(\ab[1][21] ), .IN2(\ab[0][22] ), .Q(n5) );
  AND2X1 U5 ( .IN1(\ab[1][20] ), .IN2(\ab[0][21] ), .Q(n6) );
  AND2X1 U6 ( .IN1(\ab[1][19] ), .IN2(\ab[0][20] ), .Q(n7) );
  AND2X1 U7 ( .IN1(\ab[1][18] ), .IN2(\ab[0][19] ), .Q(n8) );
  AND2X1 U8 ( .IN1(\ab[1][17] ), .IN2(\ab[0][18] ), .Q(n9) );
  AND2X1 U9 ( .IN1(\ab[1][16] ), .IN2(\ab[0][17] ), .Q(n10) );
  AND2X1 U10 ( .IN1(\ab[1][15] ), .IN2(\ab[0][16] ), .Q(n11) );
  AND2X1 U11 ( .IN1(\ab[1][14] ), .IN2(\ab[0][15] ), .Q(n12) );
  AND2X1 U12 ( .IN1(\ab[1][13] ), .IN2(\ab[0][14] ), .Q(n13) );
  AND2X1 U13 ( .IN1(\ab[1][12] ), .IN2(\ab[0][13] ), .Q(n14) );
  AND2X1 U14 ( .IN1(\ab[1][11] ), .IN2(\ab[0][12] ), .Q(n15) );
  AND2X1 U15 ( .IN1(\ab[1][10] ), .IN2(\ab[0][11] ), .Q(n16) );
  AND2X1 U16 ( .IN1(\ab[1][9] ), .IN2(\ab[0][10] ), .Q(n17) );
  AND2X1 U17 ( .IN1(\ab[1][8] ), .IN2(\ab[0][9] ), .Q(n18) );
  AND2X1 U18 ( .IN1(\ab[1][7] ), .IN2(\ab[0][8] ), .Q(n19) );
  AND2X1 U19 ( .IN1(\ab[1][6] ), .IN2(\ab[0][7] ), .Q(n20) );
  AND2X1 U20 ( .IN1(\ab[1][5] ), .IN2(\ab[0][6] ), .Q(n21) );
  AND2X1 U21 ( .IN1(\ab[1][4] ), .IN2(\ab[0][5] ), .Q(n22) );
  AND2X1 U22 ( .IN1(\ab[1][3] ), .IN2(\ab[0][4] ), .Q(n23) );
  AND2X1 U23 ( .IN1(\ab[1][2] ), .IN2(\ab[0][3] ), .Q(n24) );
  AND2X1 U24 ( .IN1(\CARRYB[23][22] ), .IN2(\ab[23][23] ), .Q(n25) );
  AND2X1 U25 ( .IN1(\CARRYB[23][21] ), .IN2(\SUMB[23][22] ), .Q(n26) );
  AND2X1 U26 ( .IN1(\CARRYB[23][10] ), .IN2(\SUMB[23][11] ), .Q(n27) );
  AND2X1 U27 ( .IN1(\CARRYB[23][11] ), .IN2(\SUMB[23][12] ), .Q(n28) );
  AND2X1 U28 ( .IN1(\CARRYB[23][12] ), .IN2(\SUMB[23][13] ), .Q(n29) );
  AND2X1 U29 ( .IN1(\CARRYB[23][13] ), .IN2(\SUMB[23][14] ), .Q(n30) );
  AND2X1 U30 ( .IN1(\CARRYB[23][14] ), .IN2(\SUMB[23][15] ), .Q(n31) );
  AND2X1 U31 ( .IN1(\CARRYB[23][15] ), .IN2(\SUMB[23][16] ), .Q(n32) );
  AND2X1 U32 ( .IN1(\CARRYB[23][16] ), .IN2(\SUMB[23][17] ), .Q(n33) );
  AND2X1 U33 ( .IN1(\CARRYB[23][17] ), .IN2(\SUMB[23][18] ), .Q(n34) );
  AND2X1 U34 ( .IN1(\CARRYB[23][18] ), .IN2(\SUMB[23][19] ), .Q(n35) );
  AND2X1 U35 ( .IN1(\CARRYB[23][19] ), .IN2(\SUMB[23][20] ), .Q(n36) );
  AND2X1 U36 ( .IN1(\CARRYB[23][20] ), .IN2(\SUMB[23][21] ), .Q(n37) );
  AND2X1 U37 ( .IN1(\CARRYB[23][2] ), .IN2(\SUMB[23][3] ), .Q(n38) );
  AND2X1 U38 ( .IN1(\CARRYB[23][3] ), .IN2(\SUMB[23][4] ), .Q(n39) );
  AND2X1 U39 ( .IN1(\CARRYB[23][4] ), .IN2(\SUMB[23][5] ), .Q(n40) );
  AND2X1 U40 ( .IN1(\CARRYB[23][5] ), .IN2(\SUMB[23][6] ), .Q(n41) );
  AND2X1 U41 ( .IN1(\CARRYB[23][6] ), .IN2(\SUMB[23][7] ), .Q(n42) );
  AND2X1 U42 ( .IN1(\CARRYB[23][7] ), .IN2(\SUMB[23][8] ), .Q(n43) );
  AND2X1 U43 ( .IN1(\CARRYB[23][8] ), .IN2(\SUMB[23][9] ), .Q(n44) );
  AND2X1 U44 ( .IN1(\CARRYB[23][9] ), .IN2(\SUMB[23][10] ), .Q(n45) );
  AND2X1 U45 ( .IN1(\CARRYB[23][1] ), .IN2(\SUMB[23][2] ), .Q(n46) );
  AND2X1 U46 ( .IN1(\CARRYB[23][0] ), .IN2(\SUMB[23][1] ), .Q(n47) );
  INVX0 U47 ( .INP(B[0]), .ZN(n116) );
  INVX0 U48 ( .INP(A[0]), .ZN(n93) );
  NBUFFX2 U49 ( .INP(n132), .Z(n83) );
  NBUFFX2 U50 ( .INP(n133), .Z(n84) );
  NBUFFX2 U51 ( .INP(n134), .Z(n85) );
  NBUFFX2 U52 ( .INP(n135), .Z(n86) );
  NBUFFX2 U53 ( .INP(n136), .Z(n87) );
  NBUFFX2 U54 ( .INP(n137), .Z(n88) );
  NBUFFX2 U55 ( .INP(n131), .Z(n82) );
  NBUFFX2 U56 ( .INP(n130), .Z(n81) );
  NBUFFX2 U57 ( .INP(n117), .Z(n69) );
  NBUFFX2 U58 ( .INP(n118), .Z(n70) );
  NBUFFX2 U59 ( .INP(n119), .Z(n71) );
  NBUFFX2 U60 ( .INP(n120), .Z(n72) );
  NBUFFX2 U61 ( .INP(n121), .Z(n73) );
  NBUFFX2 U62 ( .INP(n122), .Z(n74) );
  NBUFFX2 U63 ( .INP(n124), .Z(n76) );
  NBUFFX2 U64 ( .INP(n125), .Z(n77) );
  NBUFFX2 U65 ( .INP(n126), .Z(n78) );
  NBUFFX2 U66 ( .INP(n115), .Z(n68) );
  NBUFFX2 U67 ( .INP(n108), .Z(n61) );
  NBUFFX2 U68 ( .INP(n109), .Z(n62) );
  NBUFFX2 U69 ( .INP(n110), .Z(n63) );
  NBUFFX2 U70 ( .INP(n111), .Z(n64) );
  NBUFFX2 U71 ( .INP(n113), .Z(n66) );
  NBUFFX2 U72 ( .INP(n114), .Z(n67) );
  NBUFFX2 U73 ( .INP(n94), .Z(n48) );
  NBUFFX2 U74 ( .INP(n112), .Z(n65) );
  NBUFFX2 U75 ( .INP(n95), .Z(n49) );
  NBUFFX2 U76 ( .INP(n96), .Z(n50) );
  NBUFFX2 U77 ( .INP(n97), .Z(n51) );
  NBUFFX2 U78 ( .INP(n98), .Z(n52) );
  NBUFFX2 U79 ( .INP(n99), .Z(n53) );
  NBUFFX2 U80 ( .INP(n100), .Z(n54) );
  NBUFFX2 U81 ( .INP(n101), .Z(n55) );
  NBUFFX2 U82 ( .INP(n102), .Z(n56) );
  NBUFFX2 U83 ( .INP(n103), .Z(n57) );
  NBUFFX2 U84 ( .INP(n105), .Z(n58) );
  NBUFFX2 U85 ( .INP(n106), .Z(n59) );
  NBUFFX2 U86 ( .INP(n107), .Z(n60) );
  NBUFFX2 U87 ( .INP(n138), .Z(n89) );
  NBUFFX2 U88 ( .INP(n123), .Z(n75) );
  NBUFFX2 U89 ( .INP(n128), .Z(n79) );
  NBUFFX2 U90 ( .INP(n129), .Z(n80) );
  INVX0 U91 ( .INP(B[1]), .ZN(n127) );
  INVX0 U92 ( .INP(A[1]), .ZN(n104) );
  INVX0 U93 ( .INP(B[4]), .ZN(n133) );
  INVX0 U94 ( .INP(B[5]), .ZN(n134) );
  INVX0 U95 ( .INP(B[6]), .ZN(n135) );
  INVX0 U96 ( .INP(B[7]), .ZN(n136) );
  INVX0 U97 ( .INP(B[8]), .ZN(n137) );
  INVX0 U98 ( .INP(B[9]), .ZN(n138) );
  INVX0 U99 ( .INP(B[3]), .ZN(n132) );
  INVX0 U100 ( .INP(A[2]), .ZN(n108) );
  INVX0 U101 ( .INP(B[22]), .ZN(n130) );
  INVX0 U102 ( .INP(A[3]), .ZN(n109) );
  INVX0 U103 ( .INP(B[10]), .ZN(n117) );
  INVX0 U104 ( .INP(B[11]), .ZN(n118) );
  INVX0 U105 ( .INP(B[12]), .ZN(n119) );
  INVX0 U106 ( .INP(B[13]), .ZN(n120) );
  INVX0 U107 ( .INP(B[14]), .ZN(n121) );
  INVX0 U108 ( .INP(B[15]), .ZN(n122) );
  INVX0 U109 ( .INP(B[16]), .ZN(n123) );
  INVX0 U110 ( .INP(B[17]), .ZN(n124) );
  INVX0 U111 ( .INP(B[18]), .ZN(n125) );
  INVX0 U112 ( .INP(B[19]), .ZN(n126) );
  INVX0 U113 ( .INP(B[20]), .ZN(n128) );
  INVX0 U114 ( .INP(B[21]), .ZN(n129) );
  INVX0 U115 ( .INP(A[4]), .ZN(n110) );
  INVX0 U116 ( .INP(A[5]), .ZN(n111) );
  INVX0 U117 ( .INP(B[2]), .ZN(n131) );
  INVX0 U118 ( .INP(A[6]), .ZN(n112) );
  INVX0 U119 ( .INP(A[7]), .ZN(n113) );
  INVX0 U120 ( .INP(A[8]), .ZN(n114) );
  INVX0 U121 ( .INP(A[9]), .ZN(n115) );
  INVX0 U122 ( .INP(A[10]), .ZN(n94) );
  INVX0 U123 ( .INP(A[11]), .ZN(n95) );
  INVX0 U124 ( .INP(A[12]), .ZN(n96) );
  INVX0 U125 ( .INP(A[13]), .ZN(n97) );
  INVX0 U126 ( .INP(A[14]), .ZN(n98) );
  INVX0 U127 ( .INP(A[15]), .ZN(n99) );
  INVX0 U128 ( .INP(A[16]), .ZN(n100) );
  INVX0 U129 ( .INP(A[17]), .ZN(n101) );
  INVX0 U130 ( .INP(A[18]), .ZN(n102) );
  INVX0 U131 ( .INP(A[19]), .ZN(n103) );
  INVX0 U132 ( .INP(A[20]), .ZN(n105) );
  INVX0 U133 ( .INP(A[21]), .ZN(n106) );
  INVX0 U134 ( .INP(A[22]), .ZN(n107) );
  XOR2X1 U135 ( .IN1(\CARRYB[23][0] ), .IN2(\SUMB[23][1] ), .Q(\A1[22] ) );
  XOR2X1 U136 ( .IN1(\CARRYB[23][1] ), .IN2(\SUMB[23][2] ), .Q(\A1[23] ) );
  XOR2X1 U137 ( .IN1(\CARRYB[23][2] ), .IN2(\SUMB[23][3] ), .Q(\A1[24] ) );
  XOR2X1 U138 ( .IN1(\CARRYB[23][3] ), .IN2(\SUMB[23][4] ), .Q(\A1[25] ) );
  XOR2X1 U139 ( .IN1(\CARRYB[23][4] ), .IN2(\SUMB[23][5] ), .Q(\A1[26] ) );
  XOR2X1 U140 ( .IN1(\CARRYB[23][5] ), .IN2(\SUMB[23][6] ), .Q(\A1[27] ) );
  XOR2X1 U141 ( .IN1(\CARRYB[23][6] ), .IN2(\SUMB[23][7] ), .Q(\A1[28] ) );
  XOR2X1 U142 ( .IN1(\CARRYB[23][7] ), .IN2(\SUMB[23][8] ), .Q(\A1[29] ) );
  XOR2X1 U143 ( .IN1(\CARRYB[23][8] ), .IN2(\SUMB[23][9] ), .Q(\A1[30] ) );
  XOR2X1 U144 ( .IN1(\CARRYB[23][9] ), .IN2(\SUMB[23][10] ), .Q(\A1[31] ) );
  XOR2X1 U145 ( .IN1(\CARRYB[23][10] ), .IN2(\SUMB[23][11] ), .Q(\A1[32] ) );
  XOR2X1 U146 ( .IN1(\CARRYB[23][11] ), .IN2(\SUMB[23][12] ), .Q(\A1[33] ) );
  XOR2X1 U147 ( .IN1(\CARRYB[23][12] ), .IN2(\SUMB[23][13] ), .Q(\A1[34] ) );
  XOR2X1 U148 ( .IN1(\CARRYB[23][13] ), .IN2(\SUMB[23][14] ), .Q(\A1[35] ) );
  XOR2X1 U149 ( .IN1(\CARRYB[23][14] ), .IN2(\SUMB[23][15] ), .Q(\A1[36] ) );
  XOR2X1 U150 ( .IN1(\CARRYB[23][15] ), .IN2(\SUMB[23][16] ), .Q(\A1[37] ) );
  XOR2X1 U151 ( .IN1(\CARRYB[23][16] ), .IN2(\SUMB[23][17] ), .Q(\A1[38] ) );
  XOR2X1 U152 ( .IN1(\CARRYB[23][17] ), .IN2(\SUMB[23][18] ), .Q(\A1[39] ) );
  XOR2X1 U153 ( .IN1(\CARRYB[23][18] ), .IN2(\SUMB[23][19] ), .Q(\A1[40] ) );
  XOR2X1 U154 ( .IN1(\CARRYB[23][19] ), .IN2(\SUMB[23][20] ), .Q(\A1[41] ) );
  XOR2X1 U155 ( .IN1(\CARRYB[23][20] ), .IN2(\SUMB[23][21] ), .Q(\A1[42] ) );
  XOR2X1 U156 ( .IN1(\CARRYB[23][21] ), .IN2(\SUMB[23][22] ), .Q(\A1[43] ) );
  XOR2X1 U157 ( .IN1(\CARRYB[23][22] ), .IN2(\ab[23][23] ), .Q(\A1[44] ) );
  XOR2X1 U158 ( .IN1(\ab[0][2] ), .IN2(\ab[1][1] ), .Q(\SUMB[1][1] ) );
  XOR2X1 U159 ( .IN1(\ab[0][3] ), .IN2(\ab[1][2] ), .Q(\SUMB[1][2] ) );
  XOR2X1 U160 ( .IN1(\ab[0][4] ), .IN2(\ab[1][3] ), .Q(\SUMB[1][3] ) );
  XOR2X1 U161 ( .IN1(\ab[0][5] ), .IN2(\ab[1][4] ), .Q(\SUMB[1][4] ) );
  XOR2X1 U162 ( .IN1(\ab[0][6] ), .IN2(\ab[1][5] ), .Q(\SUMB[1][5] ) );
  XOR2X1 U163 ( .IN1(\ab[0][7] ), .IN2(\ab[1][6] ), .Q(\SUMB[1][6] ) );
  XOR2X1 U164 ( .IN1(\ab[0][8] ), .IN2(\ab[1][7] ), .Q(\SUMB[1][7] ) );
  XOR2X1 U165 ( .IN1(\ab[0][9] ), .IN2(\ab[1][8] ), .Q(\SUMB[1][8] ) );
  XOR2X1 U166 ( .IN1(\ab[0][10] ), .IN2(\ab[1][9] ), .Q(\SUMB[1][9] ) );
  XOR2X1 U167 ( .IN1(\ab[0][11] ), .IN2(\ab[1][10] ), .Q(\SUMB[1][10] ) );
  XOR2X1 U168 ( .IN1(\ab[0][12] ), .IN2(\ab[1][11] ), .Q(\SUMB[1][11] ) );
  XOR2X1 U169 ( .IN1(\ab[0][13] ), .IN2(\ab[1][12] ), .Q(\SUMB[1][12] ) );
  XOR2X1 U170 ( .IN1(\ab[0][14] ), .IN2(\ab[1][13] ), .Q(\SUMB[1][13] ) );
  XOR2X1 U171 ( .IN1(\ab[0][15] ), .IN2(\ab[1][14] ), .Q(\SUMB[1][14] ) );
  XOR2X1 U172 ( .IN1(\ab[0][16] ), .IN2(\ab[1][15] ), .Q(\SUMB[1][15] ) );
  XOR2X1 U173 ( .IN1(\ab[0][17] ), .IN2(\ab[1][16] ), .Q(\SUMB[1][16] ) );
  XOR2X1 U174 ( .IN1(\ab[0][18] ), .IN2(\ab[1][17] ), .Q(\SUMB[1][17] ) );
  XOR2X1 U175 ( .IN1(\ab[0][19] ), .IN2(\ab[1][18] ), .Q(\SUMB[1][18] ) );
  XOR2X1 U176 ( .IN1(\ab[0][20] ), .IN2(\ab[1][19] ), .Q(\SUMB[1][19] ) );
  XOR2X1 U177 ( .IN1(\ab[0][21] ), .IN2(\ab[1][20] ), .Q(\SUMB[1][20] ) );
  XOR2X1 U178 ( .IN1(\ab[0][22] ), .IN2(\ab[1][21] ), .Q(\SUMB[1][21] ) );
  XOR2X1 U179 ( .IN1(\ab[0][23] ), .IN2(\ab[1][22] ), .Q(\SUMB[1][22] ) );
  INVX0 U180 ( .INP(\ab[23][23] ), .ZN(n90) );
  INVX0 U181 ( .INP(\ab[23][23] ), .ZN(n91) );
  INVX0 U182 ( .INP(\ab[23][23] ), .ZN(n92) );
  NOR2X0 U184 ( .IN1(n68), .IN2(n138), .QN(\ab[9][9] ) );
  NOR2X0 U185 ( .IN1(n68), .IN2(n88), .QN(\ab[9][8] ) );
  NOR2X0 U186 ( .IN1(n68), .IN2(n87), .QN(\ab[9][7] ) );
  NOR2X0 U187 ( .IN1(n68), .IN2(n86), .QN(\ab[9][6] ) );
  NOR2X0 U188 ( .IN1(n68), .IN2(n85), .QN(\ab[9][5] ) );
  NOR2X0 U189 ( .IN1(n68), .IN2(n84), .QN(\ab[9][4] ) );
  NOR2X0 U190 ( .IN1(n68), .IN2(n83), .QN(\ab[9][3] ) );
  NOR2X0 U191 ( .IN1(n68), .IN2(n82), .QN(\ab[9][2] ) );
  NOR2X0 U192 ( .IN1(n68), .IN2(n90), .QN(\ab[9][23] ) );
  NOR2X0 U193 ( .IN1(n68), .IN2(n81), .QN(\ab[9][22] ) );
  NOR2X0 U194 ( .IN1(n68), .IN2(n129), .QN(\ab[9][21] ) );
  NOR2X0 U195 ( .IN1(n68), .IN2(n128), .QN(\ab[9][20] ) );
  NOR2X0 U196 ( .IN1(n115), .IN2(n127), .QN(\ab[9][1] ) );
  NOR2X0 U197 ( .IN1(n115), .IN2(n78), .QN(\ab[9][19] ) );
  NOR2X0 U198 ( .IN1(n115), .IN2(n77), .QN(\ab[9][18] ) );
  NOR2X0 U199 ( .IN1(n115), .IN2(n76), .QN(\ab[9][17] ) );
  NOR2X0 U200 ( .IN1(n115), .IN2(n123), .QN(\ab[9][16] ) );
  NOR2X0 U201 ( .IN1(n115), .IN2(n74), .QN(\ab[9][15] ) );
  NOR2X0 U202 ( .IN1(n115), .IN2(n73), .QN(\ab[9][14] ) );
  NOR2X0 U203 ( .IN1(n115), .IN2(n72), .QN(\ab[9][13] ) );
  NOR2X0 U204 ( .IN1(n115), .IN2(n71), .QN(\ab[9][12] ) );
  NOR2X0 U205 ( .IN1(n115), .IN2(n70), .QN(\ab[9][11] ) );
  NOR2X0 U206 ( .IN1(n115), .IN2(n69), .QN(\ab[9][10] ) );
  NOR2X0 U207 ( .IN1(n68), .IN2(n116), .QN(\ab[9][0] ) );
  NOR2X0 U208 ( .IN1(n89), .IN2(n67), .QN(\ab[8][9] ) );
  NOR2X0 U209 ( .IN1(n88), .IN2(n67), .QN(\ab[8][8] ) );
  NOR2X0 U210 ( .IN1(n87), .IN2(n67), .QN(\ab[8][7] ) );
  NOR2X0 U211 ( .IN1(n86), .IN2(n67), .QN(\ab[8][6] ) );
  NOR2X0 U212 ( .IN1(n85), .IN2(n67), .QN(\ab[8][5] ) );
  NOR2X0 U213 ( .IN1(n84), .IN2(n67), .QN(\ab[8][4] ) );
  NOR2X0 U214 ( .IN1(n83), .IN2(n67), .QN(\ab[8][3] ) );
  NOR2X0 U215 ( .IN1(n82), .IN2(n67), .QN(\ab[8][2] ) );
  NOR2X0 U216 ( .IN1(n91), .IN2(n67), .QN(\ab[8][23] ) );
  NOR2X0 U217 ( .IN1(n81), .IN2(n67), .QN(\ab[8][22] ) );
  NOR2X0 U218 ( .IN1(n129), .IN2(n67), .QN(\ab[8][21] ) );
  NOR2X0 U219 ( .IN1(n128), .IN2(n67), .QN(\ab[8][20] ) );
  NOR2X0 U220 ( .IN1(n127), .IN2(n114), .QN(\ab[8][1] ) );
  NOR2X0 U221 ( .IN1(n78), .IN2(n114), .QN(\ab[8][19] ) );
  NOR2X0 U222 ( .IN1(n77), .IN2(n114), .QN(\ab[8][18] ) );
  NOR2X0 U223 ( .IN1(n76), .IN2(n114), .QN(\ab[8][17] ) );
  NOR2X0 U224 ( .IN1(n123), .IN2(n114), .QN(\ab[8][16] ) );
  NOR2X0 U225 ( .IN1(n74), .IN2(n114), .QN(\ab[8][15] ) );
  NOR2X0 U226 ( .IN1(n73), .IN2(n114), .QN(\ab[8][14] ) );
  NOR2X0 U227 ( .IN1(n72), .IN2(n114), .QN(\ab[8][13] ) );
  NOR2X0 U228 ( .IN1(n71), .IN2(n114), .QN(\ab[8][12] ) );
  NOR2X0 U229 ( .IN1(n70), .IN2(n114), .QN(\ab[8][11] ) );
  NOR2X0 U230 ( .IN1(n69), .IN2(n114), .QN(\ab[8][10] ) );
  NOR2X0 U231 ( .IN1(n116), .IN2(n67), .QN(\ab[8][0] ) );
  NOR2X0 U232 ( .IN1(n138), .IN2(n66), .QN(\ab[7][9] ) );
  NOR2X0 U233 ( .IN1(n88), .IN2(n66), .QN(\ab[7][8] ) );
  NOR2X0 U234 ( .IN1(n87), .IN2(n66), .QN(\ab[7][7] ) );
  NOR2X0 U235 ( .IN1(n86), .IN2(n66), .QN(\ab[7][6] ) );
  NOR2X0 U236 ( .IN1(n85), .IN2(n66), .QN(\ab[7][5] ) );
  NOR2X0 U237 ( .IN1(n84), .IN2(n66), .QN(\ab[7][4] ) );
  NOR2X0 U238 ( .IN1(n83), .IN2(n66), .QN(\ab[7][3] ) );
  NOR2X0 U239 ( .IN1(n82), .IN2(n66), .QN(\ab[7][2] ) );
  NOR2X0 U240 ( .IN1(n92), .IN2(n66), .QN(\ab[7][23] ) );
  NOR2X0 U241 ( .IN1(n81), .IN2(n66), .QN(\ab[7][22] ) );
  NOR2X0 U242 ( .IN1(n129), .IN2(n66), .QN(\ab[7][21] ) );
  NOR2X0 U243 ( .IN1(n128), .IN2(n66), .QN(\ab[7][20] ) );
  NOR2X0 U244 ( .IN1(n127), .IN2(n113), .QN(\ab[7][1] ) );
  NOR2X0 U245 ( .IN1(n78), .IN2(n113), .QN(\ab[7][19] ) );
  NOR2X0 U246 ( .IN1(n77), .IN2(n113), .QN(\ab[7][18] ) );
  NOR2X0 U247 ( .IN1(n76), .IN2(n113), .QN(\ab[7][17] ) );
  NOR2X0 U248 ( .IN1(n123), .IN2(n113), .QN(\ab[7][16] ) );
  NOR2X0 U249 ( .IN1(n74), .IN2(n113), .QN(\ab[7][15] ) );
  NOR2X0 U250 ( .IN1(n73), .IN2(n113), .QN(\ab[7][14] ) );
  NOR2X0 U251 ( .IN1(n72), .IN2(n113), .QN(\ab[7][13] ) );
  NOR2X0 U252 ( .IN1(n71), .IN2(n113), .QN(\ab[7][12] ) );
  NOR2X0 U253 ( .IN1(n70), .IN2(n113), .QN(\ab[7][11] ) );
  NOR2X0 U254 ( .IN1(n69), .IN2(n113), .QN(\ab[7][10] ) );
  NOR2X0 U255 ( .IN1(n116), .IN2(n66), .QN(\ab[7][0] ) );
  NOR2X0 U256 ( .IN1(n89), .IN2(n112), .QN(\ab[6][9] ) );
  NOR2X0 U257 ( .IN1(n88), .IN2(n112), .QN(\ab[6][8] ) );
  NOR2X0 U258 ( .IN1(n87), .IN2(n112), .QN(\ab[6][7] ) );
  NOR2X0 U259 ( .IN1(n86), .IN2(n112), .QN(\ab[6][6] ) );
  NOR2X0 U260 ( .IN1(n85), .IN2(n112), .QN(\ab[6][5] ) );
  NOR2X0 U261 ( .IN1(n84), .IN2(n112), .QN(\ab[6][4] ) );
  NOR2X0 U262 ( .IN1(n83), .IN2(n112), .QN(\ab[6][3] ) );
  NOR2X0 U263 ( .IN1(n82), .IN2(n112), .QN(\ab[6][2] ) );
  NOR2X0 U264 ( .IN1(n91), .IN2(n112), .QN(\ab[6][23] ) );
  NOR2X0 U265 ( .IN1(n81), .IN2(n112), .QN(\ab[6][22] ) );
  NOR2X0 U266 ( .IN1(n80), .IN2(n112), .QN(\ab[6][21] ) );
  NOR2X0 U267 ( .IN1(n79), .IN2(n65), .QN(\ab[6][20] ) );
  NOR2X0 U268 ( .IN1(n127), .IN2(n65), .QN(\ab[6][1] ) );
  NOR2X0 U269 ( .IN1(n78), .IN2(n65), .QN(\ab[6][19] ) );
  NOR2X0 U270 ( .IN1(n77), .IN2(n65), .QN(\ab[6][18] ) );
  NOR2X0 U271 ( .IN1(n76), .IN2(n65), .QN(\ab[6][17] ) );
  NOR2X0 U272 ( .IN1(n75), .IN2(n65), .QN(\ab[6][16] ) );
  NOR2X0 U273 ( .IN1(n74), .IN2(n65), .QN(\ab[6][15] ) );
  NOR2X0 U274 ( .IN1(n73), .IN2(n65), .QN(\ab[6][14] ) );
  NOR2X0 U275 ( .IN1(n72), .IN2(n65), .QN(\ab[6][13] ) );
  NOR2X0 U276 ( .IN1(n71), .IN2(n65), .QN(\ab[6][12] ) );
  NOR2X0 U277 ( .IN1(n70), .IN2(n65), .QN(\ab[6][11] ) );
  NOR2X0 U278 ( .IN1(n69), .IN2(n65), .QN(\ab[6][10] ) );
  NOR2X0 U279 ( .IN1(n116), .IN2(n65), .QN(\ab[6][0] ) );
  NOR2X0 U280 ( .IN1(n138), .IN2(n64), .QN(\ab[5][9] ) );
  NOR2X0 U281 ( .IN1(n88), .IN2(n64), .QN(\ab[5][8] ) );
  NOR2X0 U282 ( .IN1(n87), .IN2(n64), .QN(\ab[5][7] ) );
  NOR2X0 U283 ( .IN1(n86), .IN2(n64), .QN(\ab[5][6] ) );
  NOR2X0 U284 ( .IN1(n85), .IN2(n64), .QN(\ab[5][5] ) );
  NOR2X0 U285 ( .IN1(n84), .IN2(n64), .QN(\ab[5][4] ) );
  NOR2X0 U286 ( .IN1(n83), .IN2(n64), .QN(\ab[5][3] ) );
  NOR2X0 U287 ( .IN1(n82), .IN2(n64), .QN(\ab[5][2] ) );
  NOR2X0 U288 ( .IN1(n90), .IN2(n64), .QN(\ab[5][23] ) );
  NOR2X0 U289 ( .IN1(n81), .IN2(n64), .QN(\ab[5][22] ) );
  NOR2X0 U290 ( .IN1(n129), .IN2(n64), .QN(\ab[5][21] ) );
  NOR2X0 U291 ( .IN1(n128), .IN2(n64), .QN(\ab[5][20] ) );
  NOR2X0 U292 ( .IN1(n127), .IN2(n111), .QN(\ab[5][1] ) );
  NOR2X0 U293 ( .IN1(n78), .IN2(n111), .QN(\ab[5][19] ) );
  NOR2X0 U294 ( .IN1(n77), .IN2(n111), .QN(\ab[5][18] ) );
  NOR2X0 U295 ( .IN1(n76), .IN2(n111), .QN(\ab[5][17] ) );
  NOR2X0 U296 ( .IN1(n123), .IN2(n111), .QN(\ab[5][16] ) );
  NOR2X0 U297 ( .IN1(n74), .IN2(n111), .QN(\ab[5][15] ) );
  NOR2X0 U298 ( .IN1(n73), .IN2(n111), .QN(\ab[5][14] ) );
  NOR2X0 U299 ( .IN1(n72), .IN2(n111), .QN(\ab[5][13] ) );
  NOR2X0 U300 ( .IN1(n71), .IN2(n111), .QN(\ab[5][12] ) );
  NOR2X0 U301 ( .IN1(n70), .IN2(n111), .QN(\ab[5][11] ) );
  NOR2X0 U302 ( .IN1(n69), .IN2(n111), .QN(\ab[5][10] ) );
  NOR2X0 U303 ( .IN1(n116), .IN2(n64), .QN(\ab[5][0] ) );
  NOR2X0 U304 ( .IN1(n138), .IN2(n63), .QN(\ab[4][9] ) );
  NOR2X0 U305 ( .IN1(n88), .IN2(n63), .QN(\ab[4][8] ) );
  NOR2X0 U306 ( .IN1(n87), .IN2(n63), .QN(\ab[4][7] ) );
  NOR2X0 U307 ( .IN1(n86), .IN2(n63), .QN(\ab[4][6] ) );
  NOR2X0 U308 ( .IN1(n85), .IN2(n63), .QN(\ab[4][5] ) );
  NOR2X0 U309 ( .IN1(n84), .IN2(n63), .QN(\ab[4][4] ) );
  NOR2X0 U310 ( .IN1(n83), .IN2(n63), .QN(\ab[4][3] ) );
  NOR2X0 U311 ( .IN1(n82), .IN2(n63), .QN(\ab[4][2] ) );
  NOR2X0 U312 ( .IN1(n92), .IN2(n63), .QN(\ab[4][23] ) );
  NOR2X0 U313 ( .IN1(n81), .IN2(n63), .QN(\ab[4][22] ) );
  NOR2X0 U314 ( .IN1(n129), .IN2(n63), .QN(\ab[4][21] ) );
  NOR2X0 U315 ( .IN1(n128), .IN2(n63), .QN(\ab[4][20] ) );
  NOR2X0 U316 ( .IN1(n127), .IN2(n110), .QN(\ab[4][1] ) );
  NOR2X0 U317 ( .IN1(n78), .IN2(n110), .QN(\ab[4][19] ) );
  NOR2X0 U318 ( .IN1(n77), .IN2(n110), .QN(\ab[4][18] ) );
  NOR2X0 U319 ( .IN1(n76), .IN2(n110), .QN(\ab[4][17] ) );
  NOR2X0 U320 ( .IN1(n123), .IN2(n110), .QN(\ab[4][16] ) );
  NOR2X0 U321 ( .IN1(n74), .IN2(n110), .QN(\ab[4][15] ) );
  NOR2X0 U322 ( .IN1(n73), .IN2(n110), .QN(\ab[4][14] ) );
  NOR2X0 U323 ( .IN1(n72), .IN2(n110), .QN(\ab[4][13] ) );
  NOR2X0 U324 ( .IN1(n71), .IN2(n110), .QN(\ab[4][12] ) );
  NOR2X0 U325 ( .IN1(n70), .IN2(n110), .QN(\ab[4][11] ) );
  NOR2X0 U326 ( .IN1(n69), .IN2(n110), .QN(\ab[4][10] ) );
  NOR2X0 U327 ( .IN1(n116), .IN2(n63), .QN(\ab[4][0] ) );
  NOR2X0 U328 ( .IN1(n138), .IN2(n62), .QN(\ab[3][9] ) );
  NOR2X0 U329 ( .IN1(n88), .IN2(n62), .QN(\ab[3][8] ) );
  NOR2X0 U330 ( .IN1(n87), .IN2(n62), .QN(\ab[3][7] ) );
  NOR2X0 U331 ( .IN1(n86), .IN2(n62), .QN(\ab[3][6] ) );
  NOR2X0 U332 ( .IN1(n85), .IN2(n62), .QN(\ab[3][5] ) );
  NOR2X0 U333 ( .IN1(n84), .IN2(n62), .QN(\ab[3][4] ) );
  NOR2X0 U334 ( .IN1(n83), .IN2(n62), .QN(\ab[3][3] ) );
  NOR2X0 U335 ( .IN1(n82), .IN2(n62), .QN(\ab[3][2] ) );
  NOR2X0 U336 ( .IN1(n91), .IN2(n62), .QN(\ab[3][23] ) );
  NOR2X0 U337 ( .IN1(n81), .IN2(n62), .QN(\ab[3][22] ) );
  NOR2X0 U338 ( .IN1(n129), .IN2(n62), .QN(\ab[3][21] ) );
  NOR2X0 U339 ( .IN1(n128), .IN2(n62), .QN(\ab[3][20] ) );
  NOR2X0 U340 ( .IN1(n127), .IN2(n109), .QN(\ab[3][1] ) );
  NOR2X0 U341 ( .IN1(n78), .IN2(n109), .QN(\ab[3][19] ) );
  NOR2X0 U342 ( .IN1(n77), .IN2(n109), .QN(\ab[3][18] ) );
  NOR2X0 U343 ( .IN1(n76), .IN2(n109), .QN(\ab[3][17] ) );
  NOR2X0 U344 ( .IN1(n123), .IN2(n109), .QN(\ab[3][16] ) );
  NOR2X0 U345 ( .IN1(n74), .IN2(n109), .QN(\ab[3][15] ) );
  NOR2X0 U346 ( .IN1(n73), .IN2(n109), .QN(\ab[3][14] ) );
  NOR2X0 U347 ( .IN1(n72), .IN2(n109), .QN(\ab[3][13] ) );
  NOR2X0 U348 ( .IN1(n71), .IN2(n109), .QN(\ab[3][12] ) );
  NOR2X0 U349 ( .IN1(n70), .IN2(n109), .QN(\ab[3][11] ) );
  NOR2X0 U350 ( .IN1(n69), .IN2(n109), .QN(\ab[3][10] ) );
  NOR2X0 U351 ( .IN1(n116), .IN2(n62), .QN(\ab[3][0] ) );
  NOR2X0 U352 ( .IN1(n138), .IN2(n61), .QN(\ab[2][9] ) );
  NOR2X0 U353 ( .IN1(n88), .IN2(n61), .QN(\ab[2][8] ) );
  NOR2X0 U354 ( .IN1(n87), .IN2(n61), .QN(\ab[2][7] ) );
  NOR2X0 U355 ( .IN1(n86), .IN2(n61), .QN(\ab[2][6] ) );
  NOR2X0 U356 ( .IN1(n85), .IN2(n61), .QN(\ab[2][5] ) );
  NOR2X0 U357 ( .IN1(n84), .IN2(n61), .QN(\ab[2][4] ) );
  NOR2X0 U358 ( .IN1(n83), .IN2(n61), .QN(\ab[2][3] ) );
  NOR2X0 U359 ( .IN1(n82), .IN2(n61), .QN(\ab[2][2] ) );
  NOR2X0 U360 ( .IN1(n90), .IN2(n61), .QN(\ab[2][23] ) );
  NOR2X0 U361 ( .IN1(n81), .IN2(n61), .QN(\ab[2][22] ) );
  NOR2X0 U362 ( .IN1(n129), .IN2(n61), .QN(\ab[2][21] ) );
  NOR2X0 U363 ( .IN1(n128), .IN2(n61), .QN(\ab[2][20] ) );
  NOR2X0 U364 ( .IN1(n127), .IN2(n108), .QN(\ab[2][1] ) );
  NOR2X0 U365 ( .IN1(n78), .IN2(n108), .QN(\ab[2][19] ) );
  NOR2X0 U366 ( .IN1(n77), .IN2(n108), .QN(\ab[2][18] ) );
  NOR2X0 U367 ( .IN1(n76), .IN2(n108), .QN(\ab[2][17] ) );
  NOR2X0 U368 ( .IN1(n123), .IN2(n108), .QN(\ab[2][16] ) );
  NOR2X0 U369 ( .IN1(n74), .IN2(n108), .QN(\ab[2][15] ) );
  NOR2X0 U370 ( .IN1(n73), .IN2(n108), .QN(\ab[2][14] ) );
  NOR2X0 U371 ( .IN1(n72), .IN2(n108), .QN(\ab[2][13] ) );
  NOR2X0 U372 ( .IN1(n71), .IN2(n108), .QN(\ab[2][12] ) );
  NOR2X0 U373 ( .IN1(n70), .IN2(n108), .QN(\ab[2][11] ) );
  NOR2X0 U374 ( .IN1(n69), .IN2(n108), .QN(\ab[2][10] ) );
  NOR2X0 U375 ( .IN1(n116), .IN2(n61), .QN(\ab[2][0] ) );
  NOR2X0 U376 ( .IN1(n138), .IN2(n90), .QN(\ab[23][9] ) );
  NOR2X0 U377 ( .IN1(n88), .IN2(n90), .QN(\ab[23][8] ) );
  NOR2X0 U378 ( .IN1(n87), .IN2(n90), .QN(\ab[23][7] ) );
  NOR2X0 U379 ( .IN1(n86), .IN2(n90), .QN(\ab[23][6] ) );
  NOR2X0 U380 ( .IN1(n85), .IN2(n90), .QN(\ab[23][5] ) );
  NOR2X0 U381 ( .IN1(n84), .IN2(n90), .QN(\ab[23][4] ) );
  NOR2X0 U382 ( .IN1(n83), .IN2(n90), .QN(\ab[23][3] ) );
  NOR2X0 U383 ( .IN1(n82), .IN2(n90), .QN(\ab[23][2] ) );
  NOR2X0 U384 ( .IN1(n92), .IN2(n81), .QN(\ab[23][22] ) );
  NOR2X0 U385 ( .IN1(n92), .IN2(n129), .QN(\ab[23][21] ) );
  NOR2X0 U386 ( .IN1(n92), .IN2(n128), .QN(\ab[23][20] ) );
  NOR2X0 U387 ( .IN1(n92), .IN2(n127), .QN(\ab[23][1] ) );
  NOR2X0 U388 ( .IN1(n92), .IN2(n78), .QN(\ab[23][19] ) );
  NOR2X0 U389 ( .IN1(n92), .IN2(n77), .QN(\ab[23][18] ) );
  NOR2X0 U390 ( .IN1(n92), .IN2(n76), .QN(\ab[23][17] ) );
  NOR2X0 U391 ( .IN1(n92), .IN2(n123), .QN(\ab[23][16] ) );
  NOR2X0 U392 ( .IN1(n92), .IN2(n74), .QN(\ab[23][15] ) );
  NOR2X0 U393 ( .IN1(n92), .IN2(n73), .QN(\ab[23][14] ) );
  NOR2X0 U394 ( .IN1(n92), .IN2(n72), .QN(\ab[23][13] ) );
  NOR2X0 U395 ( .IN1(n92), .IN2(n71), .QN(\ab[23][12] ) );
  NOR2X0 U396 ( .IN1(n92), .IN2(n70), .QN(\ab[23][11] ) );
  NOR2X0 U397 ( .IN1(n91), .IN2(n69), .QN(\ab[23][10] ) );
  NOR2X0 U398 ( .IN1(n91), .IN2(n116), .QN(\ab[23][0] ) );
  NOR2X0 U399 ( .IN1(n138), .IN2(n107), .QN(\ab[22][9] ) );
  NOR2X0 U400 ( .IN1(n88), .IN2(n107), .QN(\ab[22][8] ) );
  NOR2X0 U401 ( .IN1(n87), .IN2(n107), .QN(\ab[22][7] ) );
  NOR2X0 U402 ( .IN1(n86), .IN2(n107), .QN(\ab[22][6] ) );
  NOR2X0 U403 ( .IN1(n85), .IN2(n107), .QN(\ab[22][5] ) );
  NOR2X0 U404 ( .IN1(n84), .IN2(n107), .QN(\ab[22][4] ) );
  NOR2X0 U405 ( .IN1(n83), .IN2(n107), .QN(\ab[22][3] ) );
  NOR2X0 U406 ( .IN1(n82), .IN2(n107), .QN(\ab[22][2] ) );
  NOR2X0 U407 ( .IN1(n91), .IN2(n107), .QN(\ab[22][23] ) );
  NOR2X0 U408 ( .IN1(n81), .IN2(n107), .QN(\ab[22][22] ) );
  NOR2X0 U409 ( .IN1(n129), .IN2(n107), .QN(\ab[22][21] ) );
  NOR2X0 U410 ( .IN1(n128), .IN2(n60), .QN(\ab[22][20] ) );
  NOR2X0 U411 ( .IN1(n127), .IN2(n60), .QN(\ab[22][1] ) );
  NOR2X0 U412 ( .IN1(n78), .IN2(n60), .QN(\ab[22][19] ) );
  NOR2X0 U413 ( .IN1(n77), .IN2(n60), .QN(\ab[22][18] ) );
  NOR2X0 U414 ( .IN1(n76), .IN2(n60), .QN(\ab[22][17] ) );
  NOR2X0 U415 ( .IN1(n123), .IN2(n60), .QN(\ab[22][16] ) );
  NOR2X0 U416 ( .IN1(n74), .IN2(n60), .QN(\ab[22][15] ) );
  NOR2X0 U417 ( .IN1(n73), .IN2(n60), .QN(\ab[22][14] ) );
  NOR2X0 U418 ( .IN1(n72), .IN2(n60), .QN(\ab[22][13] ) );
  NOR2X0 U419 ( .IN1(n71), .IN2(n60), .QN(\ab[22][12] ) );
  NOR2X0 U420 ( .IN1(n70), .IN2(n60), .QN(\ab[22][11] ) );
  NOR2X0 U421 ( .IN1(n69), .IN2(n60), .QN(\ab[22][10] ) );
  NOR2X0 U422 ( .IN1(n116), .IN2(n60), .QN(\ab[22][0] ) );
  NOR2X0 U423 ( .IN1(n138), .IN2(n106), .QN(\ab[21][9] ) );
  NOR2X0 U424 ( .IN1(n88), .IN2(n106), .QN(\ab[21][8] ) );
  NOR2X0 U425 ( .IN1(n87), .IN2(n106), .QN(\ab[21][7] ) );
  NOR2X0 U426 ( .IN1(n86), .IN2(n106), .QN(\ab[21][6] ) );
  NOR2X0 U427 ( .IN1(n85), .IN2(n106), .QN(\ab[21][5] ) );
  NOR2X0 U428 ( .IN1(n84), .IN2(n106), .QN(\ab[21][4] ) );
  NOR2X0 U429 ( .IN1(n83), .IN2(n106), .QN(\ab[21][3] ) );
  NOR2X0 U430 ( .IN1(n82), .IN2(n106), .QN(\ab[21][2] ) );
  NOR2X0 U431 ( .IN1(n91), .IN2(n106), .QN(\ab[21][23] ) );
  NOR2X0 U432 ( .IN1(n81), .IN2(n106), .QN(\ab[21][22] ) );
  NOR2X0 U433 ( .IN1(n129), .IN2(n106), .QN(\ab[21][21] ) );
  NOR2X0 U434 ( .IN1(n128), .IN2(n59), .QN(\ab[21][20] ) );
  NOR2X0 U435 ( .IN1(n127), .IN2(n59), .QN(\ab[21][1] ) );
  NOR2X0 U436 ( .IN1(n78), .IN2(n59), .QN(\ab[21][19] ) );
  NOR2X0 U437 ( .IN1(n77), .IN2(n59), .QN(\ab[21][18] ) );
  NOR2X0 U438 ( .IN1(n76), .IN2(n59), .QN(\ab[21][17] ) );
  NOR2X0 U439 ( .IN1(n123), .IN2(n59), .QN(\ab[21][16] ) );
  NOR2X0 U440 ( .IN1(n74), .IN2(n59), .QN(\ab[21][15] ) );
  NOR2X0 U441 ( .IN1(n73), .IN2(n59), .QN(\ab[21][14] ) );
  NOR2X0 U442 ( .IN1(n72), .IN2(n59), .QN(\ab[21][13] ) );
  NOR2X0 U443 ( .IN1(n71), .IN2(n59), .QN(\ab[21][12] ) );
  NOR2X0 U444 ( .IN1(n70), .IN2(n59), .QN(\ab[21][11] ) );
  NOR2X0 U445 ( .IN1(n69), .IN2(n59), .QN(\ab[21][10] ) );
  NOR2X0 U446 ( .IN1(n116), .IN2(n59), .QN(\ab[21][0] ) );
  NOR2X0 U447 ( .IN1(n138), .IN2(n58), .QN(\ab[20][9] ) );
  NOR2X0 U448 ( .IN1(n88), .IN2(n58), .QN(\ab[20][8] ) );
  NOR2X0 U449 ( .IN1(n87), .IN2(n58), .QN(\ab[20][7] ) );
  NOR2X0 U450 ( .IN1(n86), .IN2(n58), .QN(\ab[20][6] ) );
  NOR2X0 U451 ( .IN1(n85), .IN2(n58), .QN(\ab[20][5] ) );
  NOR2X0 U452 ( .IN1(n84), .IN2(n58), .QN(\ab[20][4] ) );
  NOR2X0 U453 ( .IN1(n83), .IN2(n58), .QN(\ab[20][3] ) );
  NOR2X0 U454 ( .IN1(n82), .IN2(n58), .QN(\ab[20][2] ) );
  NOR2X0 U455 ( .IN1(n91), .IN2(n58), .QN(\ab[20][23] ) );
  NOR2X0 U456 ( .IN1(n81), .IN2(n58), .QN(\ab[20][22] ) );
  NOR2X0 U457 ( .IN1(n129), .IN2(n58), .QN(\ab[20][21] ) );
  NOR2X0 U458 ( .IN1(n128), .IN2(n58), .QN(\ab[20][20] ) );
  NOR2X0 U459 ( .IN1(n127), .IN2(n105), .QN(\ab[20][1] ) );
  NOR2X0 U460 ( .IN1(n78), .IN2(n105), .QN(\ab[20][19] ) );
  NOR2X0 U461 ( .IN1(n77), .IN2(n105), .QN(\ab[20][18] ) );
  NOR2X0 U462 ( .IN1(n76), .IN2(n105), .QN(\ab[20][17] ) );
  NOR2X0 U463 ( .IN1(n123), .IN2(n105), .QN(\ab[20][16] ) );
  NOR2X0 U464 ( .IN1(n74), .IN2(n105), .QN(\ab[20][15] ) );
  NOR2X0 U465 ( .IN1(n73), .IN2(n105), .QN(\ab[20][14] ) );
  NOR2X0 U466 ( .IN1(n72), .IN2(n105), .QN(\ab[20][13] ) );
  NOR2X0 U467 ( .IN1(n71), .IN2(n105), .QN(\ab[20][12] ) );
  NOR2X0 U468 ( .IN1(n70), .IN2(n105), .QN(\ab[20][11] ) );
  NOR2X0 U469 ( .IN1(n69), .IN2(n105), .QN(\ab[20][10] ) );
  NOR2X0 U470 ( .IN1(n116), .IN2(n58), .QN(\ab[20][0] ) );
  NOR2X0 U471 ( .IN1(n138), .IN2(n104), .QN(\ab[1][9] ) );
  NOR2X0 U472 ( .IN1(n88), .IN2(n104), .QN(\ab[1][8] ) );
  NOR2X0 U473 ( .IN1(n87), .IN2(n104), .QN(\ab[1][7] ) );
  NOR2X0 U474 ( .IN1(n86), .IN2(n104), .QN(\ab[1][6] ) );
  NOR2X0 U475 ( .IN1(n85), .IN2(n104), .QN(\ab[1][5] ) );
  NOR2X0 U476 ( .IN1(n84), .IN2(n104), .QN(\ab[1][4] ) );
  NOR2X0 U477 ( .IN1(n83), .IN2(n104), .QN(\ab[1][3] ) );
  NOR2X0 U478 ( .IN1(n82), .IN2(n104), .QN(\ab[1][2] ) );
  NOR2X0 U479 ( .IN1(n91), .IN2(n104), .QN(\ab[1][23] ) );
  NOR2X0 U480 ( .IN1(n130), .IN2(n104), .QN(\ab[1][22] ) );
  NOR2X0 U481 ( .IN1(n80), .IN2(n104), .QN(\ab[1][21] ) );
  NOR2X0 U482 ( .IN1(n79), .IN2(n104), .QN(\ab[1][20] ) );
  NOR2X0 U483 ( .IN1(n126), .IN2(n104), .QN(\ab[1][19] ) );
  NOR2X0 U484 ( .IN1(n125), .IN2(n104), .QN(\ab[1][18] ) );
  NOR2X0 U485 ( .IN1(n124), .IN2(n104), .QN(\ab[1][17] ) );
  NOR2X0 U486 ( .IN1(n75), .IN2(n104), .QN(\ab[1][16] ) );
  NOR2X0 U487 ( .IN1(n122), .IN2(n104), .QN(\ab[1][15] ) );
  NOR2X0 U488 ( .IN1(n121), .IN2(n104), .QN(\ab[1][14] ) );
  NOR2X0 U489 ( .IN1(n120), .IN2(n104), .QN(\ab[1][13] ) );
  NOR2X0 U490 ( .IN1(n119), .IN2(n104), .QN(\ab[1][12] ) );
  NOR2X0 U491 ( .IN1(n118), .IN2(n104), .QN(\ab[1][11] ) );
  NOR2X0 U492 ( .IN1(n117), .IN2(n104), .QN(\ab[1][10] ) );
  NOR2X0 U493 ( .IN1(n89), .IN2(n57), .QN(\ab[19][9] ) );
  NOR2X0 U494 ( .IN1(n137), .IN2(n57), .QN(\ab[19][8] ) );
  NOR2X0 U495 ( .IN1(n136), .IN2(n57), .QN(\ab[19][7] ) );
  NOR2X0 U496 ( .IN1(n135), .IN2(n57), .QN(\ab[19][6] ) );
  NOR2X0 U497 ( .IN1(n134), .IN2(n57), .QN(\ab[19][5] ) );
  NOR2X0 U498 ( .IN1(n133), .IN2(n57), .QN(\ab[19][4] ) );
  NOR2X0 U499 ( .IN1(n132), .IN2(n57), .QN(\ab[19][3] ) );
  NOR2X0 U500 ( .IN1(n131), .IN2(n57), .QN(\ab[19][2] ) );
  NOR2X0 U501 ( .IN1(n91), .IN2(n57), .QN(\ab[19][23] ) );
  NOR2X0 U502 ( .IN1(n130), .IN2(n57), .QN(\ab[19][22] ) );
  NOR2X0 U503 ( .IN1(n80), .IN2(n57), .QN(\ab[19][21] ) );
  NOR2X0 U504 ( .IN1(n79), .IN2(n57), .QN(\ab[19][20] ) );
  NOR2X0 U505 ( .IN1(n127), .IN2(n103), .QN(\ab[19][1] ) );
  NOR2X0 U506 ( .IN1(n126), .IN2(n103), .QN(\ab[19][19] ) );
  NOR2X0 U507 ( .IN1(n125), .IN2(n103), .QN(\ab[19][18] ) );
  NOR2X0 U508 ( .IN1(n124), .IN2(n103), .QN(\ab[19][17] ) );
  NOR2X0 U509 ( .IN1(n75), .IN2(n103), .QN(\ab[19][16] ) );
  NOR2X0 U510 ( .IN1(n122), .IN2(n103), .QN(\ab[19][15] ) );
  NOR2X0 U511 ( .IN1(n121), .IN2(n103), .QN(\ab[19][14] ) );
  NOR2X0 U512 ( .IN1(n120), .IN2(n103), .QN(\ab[19][13] ) );
  NOR2X0 U513 ( .IN1(n119), .IN2(n103), .QN(\ab[19][12] ) );
  NOR2X0 U514 ( .IN1(n118), .IN2(n103), .QN(\ab[19][11] ) );
  NOR2X0 U515 ( .IN1(n117), .IN2(n103), .QN(\ab[19][10] ) );
  NOR2X0 U516 ( .IN1(n116), .IN2(n57), .QN(\ab[19][0] ) );
  NOR2X0 U517 ( .IN1(n89), .IN2(n56), .QN(\ab[18][9] ) );
  NOR2X0 U518 ( .IN1(n137), .IN2(n56), .QN(\ab[18][8] ) );
  NOR2X0 U519 ( .IN1(n136), .IN2(n56), .QN(\ab[18][7] ) );
  NOR2X0 U520 ( .IN1(n135), .IN2(n56), .QN(\ab[18][6] ) );
  NOR2X0 U521 ( .IN1(n134), .IN2(n56), .QN(\ab[18][5] ) );
  NOR2X0 U522 ( .IN1(n133), .IN2(n56), .QN(\ab[18][4] ) );
  NOR2X0 U523 ( .IN1(n132), .IN2(n56), .QN(\ab[18][3] ) );
  NOR2X0 U524 ( .IN1(n131), .IN2(n56), .QN(\ab[18][2] ) );
  NOR2X0 U525 ( .IN1(n91), .IN2(n56), .QN(\ab[18][23] ) );
  NOR2X0 U526 ( .IN1(n130), .IN2(n56), .QN(\ab[18][22] ) );
  NOR2X0 U527 ( .IN1(n80), .IN2(n56), .QN(\ab[18][21] ) );
  NOR2X0 U528 ( .IN1(n79), .IN2(n56), .QN(\ab[18][20] ) );
  NOR2X0 U529 ( .IN1(n127), .IN2(n102), .QN(\ab[18][1] ) );
  NOR2X0 U530 ( .IN1(n126), .IN2(n102), .QN(\ab[18][19] ) );
  NOR2X0 U531 ( .IN1(n125), .IN2(n102), .QN(\ab[18][18] ) );
  NOR2X0 U532 ( .IN1(n124), .IN2(n102), .QN(\ab[18][17] ) );
  NOR2X0 U533 ( .IN1(n75), .IN2(n102), .QN(\ab[18][16] ) );
  NOR2X0 U534 ( .IN1(n122), .IN2(n102), .QN(\ab[18][15] ) );
  NOR2X0 U535 ( .IN1(n121), .IN2(n102), .QN(\ab[18][14] ) );
  NOR2X0 U536 ( .IN1(n120), .IN2(n102), .QN(\ab[18][13] ) );
  NOR2X0 U537 ( .IN1(n119), .IN2(n102), .QN(\ab[18][12] ) );
  NOR2X0 U538 ( .IN1(n118), .IN2(n102), .QN(\ab[18][11] ) );
  NOR2X0 U539 ( .IN1(n117), .IN2(n102), .QN(\ab[18][10] ) );
  NOR2X0 U540 ( .IN1(n116), .IN2(n56), .QN(\ab[18][0] ) );
  NOR2X0 U541 ( .IN1(n89), .IN2(n55), .QN(\ab[17][9] ) );
  NOR2X0 U542 ( .IN1(n137), .IN2(n55), .QN(\ab[17][8] ) );
  NOR2X0 U543 ( .IN1(n136), .IN2(n55), .QN(\ab[17][7] ) );
  NOR2X0 U544 ( .IN1(n135), .IN2(n55), .QN(\ab[17][6] ) );
  NOR2X0 U545 ( .IN1(n134), .IN2(n55), .QN(\ab[17][5] ) );
  NOR2X0 U546 ( .IN1(n133), .IN2(n55), .QN(\ab[17][4] ) );
  NOR2X0 U547 ( .IN1(n132), .IN2(n55), .QN(\ab[17][3] ) );
  NOR2X0 U548 ( .IN1(n131), .IN2(n55), .QN(\ab[17][2] ) );
  NOR2X0 U549 ( .IN1(n91), .IN2(n55), .QN(\ab[17][23] ) );
  NOR2X0 U550 ( .IN1(n130), .IN2(n55), .QN(\ab[17][22] ) );
  NOR2X0 U551 ( .IN1(n80), .IN2(n55), .QN(\ab[17][21] ) );
  NOR2X0 U552 ( .IN1(n79), .IN2(n55), .QN(\ab[17][20] ) );
  NOR2X0 U553 ( .IN1(n127), .IN2(n101), .QN(\ab[17][1] ) );
  NOR2X0 U554 ( .IN1(n126), .IN2(n101), .QN(\ab[17][19] ) );
  NOR2X0 U555 ( .IN1(n125), .IN2(n101), .QN(\ab[17][18] ) );
  NOR2X0 U556 ( .IN1(n124), .IN2(n101), .QN(\ab[17][17] ) );
  NOR2X0 U557 ( .IN1(n75), .IN2(n101), .QN(\ab[17][16] ) );
  NOR2X0 U558 ( .IN1(n122), .IN2(n101), .QN(\ab[17][15] ) );
  NOR2X0 U559 ( .IN1(n121), .IN2(n101), .QN(\ab[17][14] ) );
  NOR2X0 U560 ( .IN1(n120), .IN2(n101), .QN(\ab[17][13] ) );
  NOR2X0 U561 ( .IN1(n119), .IN2(n101), .QN(\ab[17][12] ) );
  NOR2X0 U562 ( .IN1(n118), .IN2(n101), .QN(\ab[17][11] ) );
  NOR2X0 U563 ( .IN1(n117), .IN2(n101), .QN(\ab[17][10] ) );
  NOR2X0 U564 ( .IN1(n116), .IN2(n55), .QN(\ab[17][0] ) );
  NOR2X0 U565 ( .IN1(n89), .IN2(n54), .QN(\ab[16][9] ) );
  NOR2X0 U566 ( .IN1(n137), .IN2(n54), .QN(\ab[16][8] ) );
  NOR2X0 U567 ( .IN1(n136), .IN2(n54), .QN(\ab[16][7] ) );
  NOR2X0 U568 ( .IN1(n135), .IN2(n54), .QN(\ab[16][6] ) );
  NOR2X0 U569 ( .IN1(n134), .IN2(n54), .QN(\ab[16][5] ) );
  NOR2X0 U570 ( .IN1(n133), .IN2(n54), .QN(\ab[16][4] ) );
  NOR2X0 U571 ( .IN1(n132), .IN2(n54), .QN(\ab[16][3] ) );
  NOR2X0 U572 ( .IN1(n131), .IN2(n54), .QN(\ab[16][2] ) );
  NOR2X0 U573 ( .IN1(n91), .IN2(n54), .QN(\ab[16][23] ) );
  NOR2X0 U574 ( .IN1(n130), .IN2(n54), .QN(\ab[16][22] ) );
  NOR2X0 U575 ( .IN1(n80), .IN2(n54), .QN(\ab[16][21] ) );
  NOR2X0 U576 ( .IN1(n79), .IN2(n54), .QN(\ab[16][20] ) );
  NOR2X0 U577 ( .IN1(n127), .IN2(n100), .QN(\ab[16][1] ) );
  NOR2X0 U578 ( .IN1(n126), .IN2(n100), .QN(\ab[16][19] ) );
  NOR2X0 U579 ( .IN1(n125), .IN2(n100), .QN(\ab[16][18] ) );
  NOR2X0 U580 ( .IN1(n124), .IN2(n100), .QN(\ab[16][17] ) );
  NOR2X0 U581 ( .IN1(n75), .IN2(n100), .QN(\ab[16][16] ) );
  NOR2X0 U582 ( .IN1(n122), .IN2(n100), .QN(\ab[16][15] ) );
  NOR2X0 U583 ( .IN1(n121), .IN2(n100), .QN(\ab[16][14] ) );
  NOR2X0 U584 ( .IN1(n120), .IN2(n100), .QN(\ab[16][13] ) );
  NOR2X0 U585 ( .IN1(n119), .IN2(n100), .QN(\ab[16][12] ) );
  NOR2X0 U586 ( .IN1(n118), .IN2(n100), .QN(\ab[16][11] ) );
  NOR2X0 U587 ( .IN1(n117), .IN2(n100), .QN(\ab[16][10] ) );
  NOR2X0 U588 ( .IN1(n116), .IN2(n54), .QN(\ab[16][0] ) );
  NOR2X0 U589 ( .IN1(n89), .IN2(n53), .QN(\ab[15][9] ) );
  NOR2X0 U590 ( .IN1(n137), .IN2(n53), .QN(\ab[15][8] ) );
  NOR2X0 U591 ( .IN1(n136), .IN2(n53), .QN(\ab[15][7] ) );
  NOR2X0 U592 ( .IN1(n135), .IN2(n53), .QN(\ab[15][6] ) );
  NOR2X0 U593 ( .IN1(n134), .IN2(n53), .QN(\ab[15][5] ) );
  NOR2X0 U594 ( .IN1(n133), .IN2(n53), .QN(\ab[15][4] ) );
  NOR2X0 U595 ( .IN1(n132), .IN2(n53), .QN(\ab[15][3] ) );
  NOR2X0 U596 ( .IN1(n131), .IN2(n53), .QN(\ab[15][2] ) );
  NOR2X0 U597 ( .IN1(n90), .IN2(n53), .QN(\ab[15][23] ) );
  NOR2X0 U598 ( .IN1(n130), .IN2(n53), .QN(\ab[15][22] ) );
  NOR2X0 U599 ( .IN1(n80), .IN2(n53), .QN(\ab[15][21] ) );
  NOR2X0 U600 ( .IN1(n79), .IN2(n53), .QN(\ab[15][20] ) );
  NOR2X0 U601 ( .IN1(n127), .IN2(n99), .QN(\ab[15][1] ) );
  NOR2X0 U602 ( .IN1(n126), .IN2(n99), .QN(\ab[15][19] ) );
  NOR2X0 U603 ( .IN1(n125), .IN2(n99), .QN(\ab[15][18] ) );
  NOR2X0 U604 ( .IN1(n124), .IN2(n99), .QN(\ab[15][17] ) );
  NOR2X0 U605 ( .IN1(n75), .IN2(n99), .QN(\ab[15][16] ) );
  NOR2X0 U606 ( .IN1(n122), .IN2(n99), .QN(\ab[15][15] ) );
  NOR2X0 U607 ( .IN1(n121), .IN2(n99), .QN(\ab[15][14] ) );
  NOR2X0 U608 ( .IN1(n120), .IN2(n99), .QN(\ab[15][13] ) );
  NOR2X0 U609 ( .IN1(n119), .IN2(n99), .QN(\ab[15][12] ) );
  NOR2X0 U610 ( .IN1(n118), .IN2(n99), .QN(\ab[15][11] ) );
  NOR2X0 U611 ( .IN1(n117), .IN2(n99), .QN(\ab[15][10] ) );
  NOR2X0 U612 ( .IN1(n116), .IN2(n53), .QN(\ab[15][0] ) );
  NOR2X0 U613 ( .IN1(n89), .IN2(n52), .QN(\ab[14][9] ) );
  NOR2X0 U614 ( .IN1(n137), .IN2(n52), .QN(\ab[14][8] ) );
  NOR2X0 U615 ( .IN1(n136), .IN2(n52), .QN(\ab[14][7] ) );
  NOR2X0 U616 ( .IN1(n135), .IN2(n52), .QN(\ab[14][6] ) );
  NOR2X0 U617 ( .IN1(n134), .IN2(n52), .QN(\ab[14][5] ) );
  NOR2X0 U618 ( .IN1(n133), .IN2(n52), .QN(\ab[14][4] ) );
  NOR2X0 U619 ( .IN1(n132), .IN2(n52), .QN(\ab[14][3] ) );
  NOR2X0 U620 ( .IN1(n131), .IN2(n52), .QN(\ab[14][2] ) );
  NOR2X0 U621 ( .IN1(n90), .IN2(n52), .QN(\ab[14][23] ) );
  NOR2X0 U622 ( .IN1(n130), .IN2(n52), .QN(\ab[14][22] ) );
  NOR2X0 U623 ( .IN1(n80), .IN2(n52), .QN(\ab[14][21] ) );
  NOR2X0 U624 ( .IN1(n79), .IN2(n52), .QN(\ab[14][20] ) );
  NOR2X0 U625 ( .IN1(n127), .IN2(n98), .QN(\ab[14][1] ) );
  NOR2X0 U626 ( .IN1(n126), .IN2(n98), .QN(\ab[14][19] ) );
  NOR2X0 U627 ( .IN1(n125), .IN2(n98), .QN(\ab[14][18] ) );
  NOR2X0 U628 ( .IN1(n124), .IN2(n98), .QN(\ab[14][17] ) );
  NOR2X0 U629 ( .IN1(n75), .IN2(n98), .QN(\ab[14][16] ) );
  NOR2X0 U630 ( .IN1(n122), .IN2(n98), .QN(\ab[14][15] ) );
  NOR2X0 U631 ( .IN1(n121), .IN2(n98), .QN(\ab[14][14] ) );
  NOR2X0 U632 ( .IN1(n120), .IN2(n98), .QN(\ab[14][13] ) );
  NOR2X0 U633 ( .IN1(n119), .IN2(n98), .QN(\ab[14][12] ) );
  NOR2X0 U634 ( .IN1(n118), .IN2(n98), .QN(\ab[14][11] ) );
  NOR2X0 U635 ( .IN1(n117), .IN2(n98), .QN(\ab[14][10] ) );
  NOR2X0 U636 ( .IN1(n116), .IN2(n52), .QN(\ab[14][0] ) );
  NOR2X0 U637 ( .IN1(n89), .IN2(n51), .QN(\ab[13][9] ) );
  NOR2X0 U638 ( .IN1(n137), .IN2(n51), .QN(\ab[13][8] ) );
  NOR2X0 U639 ( .IN1(n136), .IN2(n51), .QN(\ab[13][7] ) );
  NOR2X0 U640 ( .IN1(n135), .IN2(n51), .QN(\ab[13][6] ) );
  NOR2X0 U641 ( .IN1(n134), .IN2(n51), .QN(\ab[13][5] ) );
  NOR2X0 U642 ( .IN1(n133), .IN2(n51), .QN(\ab[13][4] ) );
  NOR2X0 U643 ( .IN1(n132), .IN2(n51), .QN(\ab[13][3] ) );
  NOR2X0 U644 ( .IN1(n131), .IN2(n51), .QN(\ab[13][2] ) );
  NOR2X0 U645 ( .IN1(n90), .IN2(n51), .QN(\ab[13][23] ) );
  NOR2X0 U646 ( .IN1(n130), .IN2(n51), .QN(\ab[13][22] ) );
  NOR2X0 U647 ( .IN1(n80), .IN2(n51), .QN(\ab[13][21] ) );
  NOR2X0 U648 ( .IN1(n79), .IN2(n51), .QN(\ab[13][20] ) );
  NOR2X0 U649 ( .IN1(n127), .IN2(n97), .QN(\ab[13][1] ) );
  NOR2X0 U650 ( .IN1(n126), .IN2(n97), .QN(\ab[13][19] ) );
  NOR2X0 U651 ( .IN1(n125), .IN2(n97), .QN(\ab[13][18] ) );
  NOR2X0 U652 ( .IN1(n124), .IN2(n97), .QN(\ab[13][17] ) );
  NOR2X0 U653 ( .IN1(n75), .IN2(n97), .QN(\ab[13][16] ) );
  NOR2X0 U654 ( .IN1(n122), .IN2(n97), .QN(\ab[13][15] ) );
  NOR2X0 U655 ( .IN1(n121), .IN2(n97), .QN(\ab[13][14] ) );
  NOR2X0 U656 ( .IN1(n120), .IN2(n97), .QN(\ab[13][13] ) );
  NOR2X0 U657 ( .IN1(n119), .IN2(n97), .QN(\ab[13][12] ) );
  NOR2X0 U658 ( .IN1(n118), .IN2(n97), .QN(\ab[13][11] ) );
  NOR2X0 U659 ( .IN1(n117), .IN2(n97), .QN(\ab[13][10] ) );
  NOR2X0 U660 ( .IN1(n116), .IN2(n51), .QN(\ab[13][0] ) );
  NOR2X0 U661 ( .IN1(n89), .IN2(n50), .QN(\ab[12][9] ) );
  NOR2X0 U662 ( .IN1(n137), .IN2(n50), .QN(\ab[12][8] ) );
  NOR2X0 U663 ( .IN1(n136), .IN2(n50), .QN(\ab[12][7] ) );
  NOR2X0 U664 ( .IN1(n135), .IN2(n50), .QN(\ab[12][6] ) );
  NOR2X0 U665 ( .IN1(n134), .IN2(n50), .QN(\ab[12][5] ) );
  NOR2X0 U666 ( .IN1(n133), .IN2(n50), .QN(\ab[12][4] ) );
  NOR2X0 U667 ( .IN1(n132), .IN2(n50), .QN(\ab[12][3] ) );
  NOR2X0 U668 ( .IN1(n131), .IN2(n50), .QN(\ab[12][2] ) );
  NOR2X0 U669 ( .IN1(n91), .IN2(n50), .QN(\ab[12][23] ) );
  NOR2X0 U670 ( .IN1(n130), .IN2(n50), .QN(\ab[12][22] ) );
  NOR2X0 U671 ( .IN1(n80), .IN2(n50), .QN(\ab[12][21] ) );
  NOR2X0 U672 ( .IN1(n79), .IN2(n50), .QN(\ab[12][20] ) );
  NOR2X0 U673 ( .IN1(n127), .IN2(n96), .QN(\ab[12][1] ) );
  NOR2X0 U674 ( .IN1(n126), .IN2(n96), .QN(\ab[12][19] ) );
  NOR2X0 U675 ( .IN1(n125), .IN2(n96), .QN(\ab[12][18] ) );
  NOR2X0 U676 ( .IN1(n124), .IN2(n96), .QN(\ab[12][17] ) );
  NOR2X0 U677 ( .IN1(n75), .IN2(n96), .QN(\ab[12][16] ) );
  NOR2X0 U678 ( .IN1(n122), .IN2(n96), .QN(\ab[12][15] ) );
  NOR2X0 U679 ( .IN1(n121), .IN2(n96), .QN(\ab[12][14] ) );
  NOR2X0 U680 ( .IN1(n120), .IN2(n96), .QN(\ab[12][13] ) );
  NOR2X0 U681 ( .IN1(n119), .IN2(n96), .QN(\ab[12][12] ) );
  NOR2X0 U682 ( .IN1(n118), .IN2(n96), .QN(\ab[12][11] ) );
  NOR2X0 U683 ( .IN1(n117), .IN2(n96), .QN(\ab[12][10] ) );
  NOR2X0 U684 ( .IN1(n116), .IN2(n50), .QN(\ab[12][0] ) );
  NOR2X0 U685 ( .IN1(n89), .IN2(n49), .QN(\ab[11][9] ) );
  NOR2X0 U686 ( .IN1(n137), .IN2(n49), .QN(\ab[11][8] ) );
  NOR2X0 U687 ( .IN1(n136), .IN2(n49), .QN(\ab[11][7] ) );
  NOR2X0 U688 ( .IN1(n135), .IN2(n49), .QN(\ab[11][6] ) );
  NOR2X0 U689 ( .IN1(n134), .IN2(n49), .QN(\ab[11][5] ) );
  NOR2X0 U690 ( .IN1(n133), .IN2(n49), .QN(\ab[11][4] ) );
  NOR2X0 U691 ( .IN1(n132), .IN2(n49), .QN(\ab[11][3] ) );
  NOR2X0 U692 ( .IN1(n131), .IN2(n49), .QN(\ab[11][2] ) );
  NOR2X0 U693 ( .IN1(n90), .IN2(n49), .QN(\ab[11][23] ) );
  NOR2X0 U694 ( .IN1(n130), .IN2(n49), .QN(\ab[11][22] ) );
  NOR2X0 U695 ( .IN1(n80), .IN2(n49), .QN(\ab[11][21] ) );
  NOR2X0 U696 ( .IN1(n79), .IN2(n49), .QN(\ab[11][20] ) );
  NOR2X0 U697 ( .IN1(n127), .IN2(n95), .QN(\ab[11][1] ) );
  NOR2X0 U698 ( .IN1(n126), .IN2(n95), .QN(\ab[11][19] ) );
  NOR2X0 U699 ( .IN1(n125), .IN2(n95), .QN(\ab[11][18] ) );
  NOR2X0 U700 ( .IN1(n124), .IN2(n95), .QN(\ab[11][17] ) );
  NOR2X0 U701 ( .IN1(n75), .IN2(n95), .QN(\ab[11][16] ) );
  NOR2X0 U702 ( .IN1(n122), .IN2(n95), .QN(\ab[11][15] ) );
  NOR2X0 U703 ( .IN1(n121), .IN2(n95), .QN(\ab[11][14] ) );
  NOR2X0 U704 ( .IN1(n120), .IN2(n95), .QN(\ab[11][13] ) );
  NOR2X0 U705 ( .IN1(n119), .IN2(n95), .QN(\ab[11][12] ) );
  NOR2X0 U706 ( .IN1(n118), .IN2(n95), .QN(\ab[11][11] ) );
  NOR2X0 U707 ( .IN1(n117), .IN2(n95), .QN(\ab[11][10] ) );
  NOR2X0 U708 ( .IN1(n116), .IN2(n49), .QN(\ab[11][0] ) );
  NOR2X0 U709 ( .IN1(n89), .IN2(n48), .QN(\ab[10][9] ) );
  NOR2X0 U710 ( .IN1(n137), .IN2(n48), .QN(\ab[10][8] ) );
  NOR2X0 U711 ( .IN1(n136), .IN2(n48), .QN(\ab[10][7] ) );
  NOR2X0 U712 ( .IN1(n135), .IN2(n48), .QN(\ab[10][6] ) );
  NOR2X0 U713 ( .IN1(n134), .IN2(n48), .QN(\ab[10][5] ) );
  NOR2X0 U714 ( .IN1(n133), .IN2(n48), .QN(\ab[10][4] ) );
  NOR2X0 U715 ( .IN1(n132), .IN2(n48), .QN(\ab[10][3] ) );
  NOR2X0 U716 ( .IN1(n131), .IN2(n48), .QN(\ab[10][2] ) );
  NOR2X0 U717 ( .IN1(n91), .IN2(n48), .QN(\ab[10][23] ) );
  NOR2X0 U718 ( .IN1(n130), .IN2(n48), .QN(\ab[10][22] ) );
  NOR2X0 U719 ( .IN1(n80), .IN2(n48), .QN(\ab[10][21] ) );
  NOR2X0 U720 ( .IN1(n79), .IN2(n48), .QN(\ab[10][20] ) );
  NOR2X0 U721 ( .IN1(n127), .IN2(n94), .QN(\ab[10][1] ) );
  NOR2X0 U722 ( .IN1(n126), .IN2(n94), .QN(\ab[10][19] ) );
  NOR2X0 U723 ( .IN1(n125), .IN2(n94), .QN(\ab[10][18] ) );
  NOR2X0 U724 ( .IN1(n124), .IN2(n94), .QN(\ab[10][17] ) );
  NOR2X0 U725 ( .IN1(n75), .IN2(n94), .QN(\ab[10][16] ) );
  NOR2X0 U726 ( .IN1(n122), .IN2(n94), .QN(\ab[10][15] ) );
  NOR2X0 U727 ( .IN1(n121), .IN2(n94), .QN(\ab[10][14] ) );
  NOR2X0 U728 ( .IN1(n120), .IN2(n94), .QN(\ab[10][13] ) );
  NOR2X0 U729 ( .IN1(n119), .IN2(n94), .QN(\ab[10][12] ) );
  NOR2X0 U730 ( .IN1(n118), .IN2(n94), .QN(\ab[10][11] ) );
  NOR2X0 U731 ( .IN1(n117), .IN2(n94), .QN(\ab[10][10] ) );
  NOR2X0 U732 ( .IN1(n116), .IN2(n48), .QN(\ab[10][0] ) );
  NOR2X0 U733 ( .IN1(n89), .IN2(n93), .QN(\ab[0][9] ) );
  NOR2X0 U734 ( .IN1(n137), .IN2(n93), .QN(\ab[0][8] ) );
  NOR2X0 U735 ( .IN1(n136), .IN2(n93), .QN(\ab[0][7] ) );
  NOR2X0 U736 ( .IN1(n135), .IN2(n93), .QN(\ab[0][6] ) );
  NOR2X0 U737 ( .IN1(n134), .IN2(n93), .QN(\ab[0][5] ) );
  NOR2X0 U738 ( .IN1(n133), .IN2(n93), .QN(\ab[0][4] ) );
  NOR2X0 U739 ( .IN1(n132), .IN2(n93), .QN(\ab[0][3] ) );
  NOR2X0 U740 ( .IN1(n131), .IN2(n93), .QN(\ab[0][2] ) );
  NOR2X0 U741 ( .IN1(n92), .IN2(n93), .QN(\ab[0][23] ) );
  NOR2X0 U742 ( .IN1(n81), .IN2(n93), .QN(\ab[0][22] ) );
  NOR2X0 U743 ( .IN1(n80), .IN2(n93), .QN(\ab[0][21] ) );
  NOR2X0 U744 ( .IN1(n79), .IN2(n93), .QN(\ab[0][20] ) );
  NOR2X0 U745 ( .IN1(n78), .IN2(n93), .QN(\ab[0][19] ) );
  NOR2X0 U746 ( .IN1(n77), .IN2(n93), .QN(\ab[0][18] ) );
  NOR2X0 U747 ( .IN1(n76), .IN2(n93), .QN(\ab[0][17] ) );
  NOR2X0 U748 ( .IN1(n75), .IN2(n93), .QN(\ab[0][16] ) );
  NOR2X0 U749 ( .IN1(n74), .IN2(n93), .QN(\ab[0][15] ) );
  NOR2X0 U750 ( .IN1(n73), .IN2(n93), .QN(\ab[0][14] ) );
  NOR2X0 U751 ( .IN1(n72), .IN2(n93), .QN(\ab[0][13] ) );
  NOR2X0 U752 ( .IN1(n71), .IN2(n93), .QN(\ab[0][12] ) );
  NOR2X0 U753 ( .IN1(n70), .IN2(n93), .QN(\ab[0][11] ) );
  NOR2X0 U754 ( .IN1(n69), .IN2(n93), .QN(\ab[0][10] ) );
  AND3X1 U755 ( .IN1(\ab[1][1] ), .IN2(B[0]), .IN3(A[0]), .Q(\CARRYB[1][0] )
         );
  NOR2X0 U756 ( .IN1(n104), .IN2(n127), .QN(\ab[1][1] ) );
endmodule


module fpalu_multiplier_DW01_inc_2 ( A, SUM );
  input [24:0] A;
  output [24:0] SUM;

  wire   [24:2] carry;

  HADDX1 U1_1_23 ( .A0(A[23]), .B0(carry[23]), .C1(SUM[24]), .SO(SUM[23]) );
  HADDX1 U1_1_22 ( .A0(A[22]), .B0(carry[22]), .C1(carry[23]), .SO(SUM[22]) );
  HADDX1 U1_1_21 ( .A0(A[21]), .B0(carry[21]), .C1(carry[22]), .SO(SUM[21]) );
  HADDX1 U1_1_20 ( .A0(A[20]), .B0(carry[20]), .C1(carry[21]), .SO(SUM[20]) );
  HADDX1 U1_1_19 ( .A0(A[19]), .B0(carry[19]), .C1(carry[20]), .SO(SUM[19]) );
  HADDX1 U1_1_18 ( .A0(A[18]), .B0(carry[18]), .C1(carry[19]), .SO(SUM[18]) );
  HADDX1 U1_1_17 ( .A0(A[17]), .B0(carry[17]), .C1(carry[18]), .SO(SUM[17]) );
  HADDX1 U1_1_16 ( .A0(A[16]), .B0(carry[16]), .C1(carry[17]), .SO(SUM[16]) );
  HADDX1 U1_1_15 ( .A0(A[15]), .B0(carry[15]), .C1(carry[16]), .SO(SUM[15]) );
  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
endmodule


module fpalu_multiplier_DW01_add_0 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [8:1] carry;

  FADDX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  FADDX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FADDX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  FADDX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X1 U1 ( .IN1(A[0]), .IN2(B[0]), .Q(n1) );
  XOR2X1 U2 ( .IN1(B[8]), .IN2(carry[8]), .Q(SUM[8]) );
  XOR2X1 U3 ( .IN1(A[0]), .IN2(B[0]), .Q(SUM[0]) );
endmodule


module fpalu_multiplier ( Ain, Bin, product, flag );
  input [31:0] Ain;
  input [31:0] Bin;
  output [31:0] product;
  output flag;
  wire   N17, N18, N19, N20, N21, N22, N23, N24, N25, N33, N34, N35, N36, N37,
         N38, N39, N40, N41, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54,
         N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68,
         N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82,
         N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N97, N98,
         N99, N100, N101, N102, N103, N104, N105, N9, N8, N15, N14, N13, N12,
         N11, N10, \sub_1_root_sub_0_root_sub_19/carry[2] ,
         \sub_1_root_sub_0_root_sub_19/carry[3] ,
         \sub_1_root_sub_0_root_sub_19/carry[4] ,
         \sub_1_root_sub_0_root_sub_19/carry[5] ,
         \sub_1_root_sub_0_root_sub_19/carry[6] ,
         \sub_1_root_sub_0_root_sub_19/carry[7] , n1, n2, n3, n4, n5, n6, n7,
         n8, n10, n11, n12, n13, n14, n15;
  wire   [8:0] exp;
  wire   [22:0] a;
  wire   [23:0] b;
  wire   [47:23] s;
  wire   [8:0] fexp1;
  wire   [24:0] sum1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22;

  LATCHX1 \sum1_reg[24]  ( .CLK(s[47]), .D(N94), .Q(sum1[24]) );
  LATCHX1 \sum1_reg[23]  ( .CLK(s[47]), .D(N93), .Q(sum1[23]) );
  LATCHX1 \sum1_reg[22]  ( .CLK(s[47]), .D(N92), .Q(sum1[22]) );
  LATCHX1 \sum1_reg[21]  ( .CLK(s[47]), .D(N91), .Q(sum1[21]) );
  LATCHX1 \sum1_reg[20]  ( .CLK(s[47]), .D(N90), .Q(sum1[20]) );
  LATCHX1 \sum1_reg[19]  ( .CLK(s[47]), .D(N89), .Q(sum1[19]) );
  LATCHX1 \sum1_reg[18]  ( .CLK(s[47]), .D(N88), .Q(sum1[18]) );
  LATCHX1 \sum1_reg[17]  ( .CLK(s[47]), .D(N87), .Q(sum1[17]) );
  LATCHX1 \sum1_reg[16]  ( .CLK(s[47]), .D(N86), .Q(sum1[16]) );
  LATCHX1 \sum1_reg[15]  ( .CLK(s[47]), .D(N85), .Q(sum1[15]) );
  LATCHX1 \sum1_reg[14]  ( .CLK(s[47]), .D(N84), .Q(sum1[14]) );
  LATCHX1 \sum1_reg[13]  ( .CLK(s[47]), .D(N83), .Q(sum1[13]) );
  LATCHX1 \sum1_reg[12]  ( .CLK(s[47]), .D(N82), .Q(sum1[12]) );
  LATCHX1 \sum1_reg[11]  ( .CLK(s[47]), .D(N81), .Q(sum1[11]) );
  LATCHX1 \sum1_reg[10]  ( .CLK(s[47]), .D(N80), .Q(sum1[10]) );
  LATCHX1 \sum1_reg[9]  ( .CLK(s[47]), .D(N79), .Q(sum1[9]) );
  LATCHX1 \sum1_reg[8]  ( .CLK(s[47]), .D(N78), .Q(sum1[8]) );
  LATCHX1 \sum1_reg[7]  ( .CLK(s[47]), .D(N77), .Q(sum1[7]) );
  LATCHX1 \sum1_reg[6]  ( .CLK(s[47]), .D(N76), .Q(sum1[6]) );
  LATCHX1 \sum1_reg[5]  ( .CLK(s[47]), .D(N75), .Q(sum1[5]) );
  LATCHX1 \sum1_reg[4]  ( .CLK(s[47]), .D(N74), .Q(sum1[4]) );
  LATCHX1 \sum1_reg[3]  ( .CLK(s[47]), .D(N73), .Q(sum1[3]) );
  LATCHX1 \sum1_reg[2]  ( .CLK(s[47]), .D(N72), .Q(sum1[2]) );
  LATCHX1 \sum1_reg[1]  ( .CLK(s[47]), .D(N71), .Q(sum1[1]) );
  LATCHX1 \sum1_reg[0]  ( .CLK(s[47]), .D(N70), .Q(sum1[0]) );
  fpalu_multiplier_DW01_inc_0 add_73 ( .A(fexp1), .SUM({N105, N104, N103, N102, 
        N101, N100, N99, N98, N97}) );
  fpalu_multiplier_DW01_inc_1 add_43 ( .A({1'b0, exp[7:0]}), .SUM({N41, N40, 
        N39, N38, N37, N36, N35, N34, N33}) );
  fpalu_multiplier_DW02_mult_0 mult_37 ( .A({n3, a}), .B({n4, b[22:0]}), .TC(
        1'b0), .PRODUCT({s, SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22}) );
  fpalu_multiplier_DW01_inc_2 add_54 ( .A({1'b0, s[47:24]}), .SUM({N69, N68, 
        N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, 
        N53, N52, N51, N50, N49, N48, N47, N46, N45}) );
  fpalu_multiplier_DW01_add_0 add_0_root_sub_0_root_sub_19 ( .A({1'b0, 
        Bin[30:23]}), .B({n2, N15, N14, N13, N12, N11, N10, N9, N8}), .CI(1'b0), .SUM({N25, N24, N23, N22, N21, N20, N19, N18, N17}) );
  MUX21X1 U3 ( .IN1(sum1[22]), .IN2(sum1[23]), .S(sum1[24]), .Q(product[22])
         );
  INVX0 U4 ( .INP(s[47]), .ZN(n8) );
  NBUFFX2 U5 ( .INP(s[23]), .Z(n7) );
  NBUFFX8 U6 ( .INP(n4), .Z(n3) );
  INVX0 U7 ( .INP(n1), .ZN(n4) );
  OR2X1 U8 ( .IN1(N25), .IN2(n11), .Q(n1) );
  NBUFFX2 U9 ( .INP(sum1[24]), .Z(n6) );
  NBUFFX2 U10 ( .INP(sum1[24]), .Z(n5) );
  INVX0 U11 ( .INP(Ain[23]), .ZN(N8) );
  NOR2X0 U12 ( .IN1(Ain[30]), .IN2(\sub_1_root_sub_0_root_sub_19/carry[7] ), 
        .QN(n2) );
  XNOR2X1 U13 ( .IN1(\sub_1_root_sub_0_root_sub_19/carry[7] ), .IN2(Ain[30]), 
        .Q(N15) );
  AND2X1 U14 ( .IN1(\sub_1_root_sub_0_root_sub_19/carry[6] ), .IN2(Ain[29]), 
        .Q(\sub_1_root_sub_0_root_sub_19/carry[7] ) );
  XOR2X1 U15 ( .IN1(Ain[29]), .IN2(\sub_1_root_sub_0_root_sub_19/carry[6] ), 
        .Q(N14) );
  AND2X1 U16 ( .IN1(\sub_1_root_sub_0_root_sub_19/carry[5] ), .IN2(Ain[28]), 
        .Q(\sub_1_root_sub_0_root_sub_19/carry[6] ) );
  XOR2X1 U17 ( .IN1(Ain[28]), .IN2(\sub_1_root_sub_0_root_sub_19/carry[5] ), 
        .Q(N13) );
  AND2X1 U18 ( .IN1(\sub_1_root_sub_0_root_sub_19/carry[4] ), .IN2(Ain[27]), 
        .Q(\sub_1_root_sub_0_root_sub_19/carry[5] ) );
  XOR2X1 U19 ( .IN1(Ain[27]), .IN2(\sub_1_root_sub_0_root_sub_19/carry[4] ), 
        .Q(N12) );
  AND2X1 U20 ( .IN1(\sub_1_root_sub_0_root_sub_19/carry[3] ), .IN2(Ain[26]), 
        .Q(\sub_1_root_sub_0_root_sub_19/carry[4] ) );
  XOR2X1 U21 ( .IN1(Ain[26]), .IN2(\sub_1_root_sub_0_root_sub_19/carry[3] ), 
        .Q(N11) );
  AND2X1 U22 ( .IN1(\sub_1_root_sub_0_root_sub_19/carry[2] ), .IN2(Ain[25]), 
        .Q(\sub_1_root_sub_0_root_sub_19/carry[3] ) );
  XOR2X1 U23 ( .IN1(Ain[25]), .IN2(\sub_1_root_sub_0_root_sub_19/carry[2] ), 
        .Q(N10) );
  AND2X1 U24 ( .IN1(Ain[23]), .IN2(Ain[24]), .Q(
        \sub_1_root_sub_0_root_sub_19/carry[2] ) );
  XOR2X1 U25 ( .IN1(Ain[24]), .IN2(Ain[23]), .Q(N9) );
  MUX21X1 U26 ( .IN1(sum1[9]), .IN2(sum1[10]), .S(n5), .Q(product[9]) );
  MUX21X1 U27 ( .IN1(sum1[8]), .IN2(sum1[9]), .S(n5), .Q(product[8]) );
  MUX21X1 U28 ( .IN1(sum1[7]), .IN2(sum1[8]), .S(n5), .Q(product[7]) );
  MUX21X1 U29 ( .IN1(sum1[6]), .IN2(sum1[7]), .S(n5), .Q(product[6]) );
  MUX21X1 U30 ( .IN1(sum1[5]), .IN2(sum1[6]), .S(n5), .Q(product[5]) );
  MUX21X1 U31 ( .IN1(sum1[4]), .IN2(sum1[5]), .S(n5), .Q(product[4]) );
  MUX21X1 U32 ( .IN1(sum1[3]), .IN2(sum1[4]), .S(n5), .Q(product[3]) );
  NOR2X0 U33 ( .IN1(n10), .IN2(n1), .QN(product[31]) );
  XNOR2X1 U34 ( .IN1(Bin[31]), .IN2(Ain[31]), .Q(n10) );
  MUX21X1 U35 ( .IN1(fexp1[7]), .IN2(N104), .S(n5), .Q(product[30]) );
  MUX21X1 U36 ( .IN1(sum1[2]), .IN2(sum1[3]), .S(n5), .Q(product[2]) );
  MUX21X1 U37 ( .IN1(fexp1[6]), .IN2(N103), .S(n5), .Q(product[29]) );
  MUX21X1 U38 ( .IN1(fexp1[5]), .IN2(N102), .S(n5), .Q(product[28]) );
  MUX21X1 U39 ( .IN1(fexp1[4]), .IN2(N101), .S(n5), .Q(product[27]) );
  MUX21X1 U40 ( .IN1(fexp1[3]), .IN2(N100), .S(n6), .Q(product[26]) );
  MUX21X1 U41 ( .IN1(fexp1[2]), .IN2(N99), .S(n6), .Q(product[25]) );
  MUX21X1 U42 ( .IN1(fexp1[1]), .IN2(N98), .S(n6), .Q(product[24]) );
  MUX21X1 U43 ( .IN1(fexp1[0]), .IN2(N97), .S(n6), .Q(product[23]) );
  MUX21X1 U44 ( .IN1(sum1[21]), .IN2(sum1[22]), .S(n6), .Q(product[21]) );
  MUX21X1 U45 ( .IN1(sum1[20]), .IN2(sum1[21]), .S(n6), .Q(product[20]) );
  MUX21X1 U46 ( .IN1(sum1[1]), .IN2(sum1[2]), .S(n6), .Q(product[1]) );
  MUX21X1 U47 ( .IN1(sum1[19]), .IN2(sum1[20]), .S(n6), .Q(product[19]) );
  MUX21X1 U48 ( .IN1(sum1[18]), .IN2(sum1[19]), .S(n6), .Q(product[18]) );
  MUX21X1 U49 ( .IN1(sum1[17]), .IN2(sum1[18]), .S(n6), .Q(product[17]) );
  MUX21X1 U50 ( .IN1(sum1[16]), .IN2(sum1[17]), .S(n6), .Q(product[16]) );
  MUX21X1 U51 ( .IN1(sum1[15]), .IN2(sum1[16]), .S(sum1[24]), .Q(product[15])
         );
  MUX21X1 U52 ( .IN1(sum1[14]), .IN2(sum1[15]), .S(sum1[24]), .Q(product[14])
         );
  MUX21X1 U53 ( .IN1(sum1[13]), .IN2(sum1[14]), .S(sum1[24]), .Q(product[13])
         );
  MUX21X1 U54 ( .IN1(sum1[12]), .IN2(sum1[13]), .S(sum1[24]), .Q(product[12])
         );
  MUX21X1 U55 ( .IN1(sum1[11]), .IN2(sum1[12]), .S(sum1[24]), .Q(product[11])
         );
  MUX21X1 U56 ( .IN1(sum1[10]), .IN2(sum1[11]), .S(sum1[24]), .Q(product[10])
         );
  MUX21X1 U57 ( .IN1(sum1[0]), .IN2(sum1[1]), .S(sum1[24]), .Q(product[0]) );
  AO221X1 U58 ( .IN1(N41), .IN2(s[47]), .IN3(N105), .IN4(sum1[24]), .IN5(n1), 
        .Q(flag) );
  AND2X1 U59 ( .IN1(s[47]), .IN2(N41), .Q(fexp1[8]) );
  MUX21X1 U60 ( .IN1(N40), .IN2(exp[7]), .S(n8), .Q(fexp1[7]) );
  MUX21X1 U61 ( .IN1(N39), .IN2(exp[6]), .S(n8), .Q(fexp1[6]) );
  MUX21X1 U62 ( .IN1(N38), .IN2(exp[5]), .S(n8), .Q(fexp1[5]) );
  MUX21X1 U63 ( .IN1(N37), .IN2(exp[4]), .S(n8), .Q(fexp1[4]) );
  MUX21X1 U64 ( .IN1(N36), .IN2(exp[3]), .S(n8), .Q(fexp1[3]) );
  MUX21X1 U65 ( .IN1(N35), .IN2(exp[2]), .S(n8), .Q(fexp1[2]) );
  MUX21X1 U66 ( .IN1(exp[1]), .IN2(N34), .S(s[47]), .Q(fexp1[1]) );
  MUX21X1 U67 ( .IN1(exp[0]), .IN2(N33), .S(s[47]), .Q(fexp1[0]) );
  AND2X1 U69 ( .IN1(n3), .IN2(N24), .Q(exp[7]) );
  AND2X1 U70 ( .IN1(n3), .IN2(N23), .Q(exp[6]) );
  AND2X1 U71 ( .IN1(n3), .IN2(N22), .Q(exp[5]) );
  AND2X1 U72 ( .IN1(n3), .IN2(N21), .Q(exp[4]) );
  AND2X1 U73 ( .IN1(n3), .IN2(N20), .Q(exp[3]) );
  AND2X1 U74 ( .IN1(n3), .IN2(N19), .Q(exp[2]) );
  AND2X1 U75 ( .IN1(n3), .IN2(N18), .Q(exp[1]) );
  AND2X1 U76 ( .IN1(n3), .IN2(N17), .Q(exp[0]) );
  AND2X1 U77 ( .IN1(Bin[9]), .IN2(n3), .Q(b[9]) );
  AND2X1 U78 ( .IN1(Bin[8]), .IN2(n3), .Q(b[8]) );
  AND2X1 U79 ( .IN1(Bin[7]), .IN2(n3), .Q(b[7]) );
  AND2X1 U80 ( .IN1(Bin[6]), .IN2(n3), .Q(b[6]) );
  AND2X1 U81 ( .IN1(Bin[5]), .IN2(n3), .Q(b[5]) );
  AND2X1 U82 ( .IN1(Bin[4]), .IN2(n3), .Q(b[4]) );
  AND2X1 U83 ( .IN1(Bin[3]), .IN2(n3), .Q(b[3]) );
  AND2X1 U84 ( .IN1(Bin[2]), .IN2(n3), .Q(b[2]) );
  AND2X1 U85 ( .IN1(Bin[22]), .IN2(n3), .Q(b[22]) );
  AND2X1 U86 ( .IN1(Bin[21]), .IN2(n3), .Q(b[21]) );
  AND2X1 U87 ( .IN1(Bin[20]), .IN2(n3), .Q(b[20]) );
  AND2X1 U88 ( .IN1(Bin[1]), .IN2(n3), .Q(b[1]) );
  AND2X1 U89 ( .IN1(Bin[19]), .IN2(n3), .Q(b[19]) );
  AND2X1 U90 ( .IN1(Bin[18]), .IN2(n3), .Q(b[18]) );
  AND2X1 U91 ( .IN1(Bin[17]), .IN2(n3), .Q(b[17]) );
  AND2X1 U92 ( .IN1(Bin[16]), .IN2(n3), .Q(b[16]) );
  AND2X1 U93 ( .IN1(Bin[15]), .IN2(n3), .Q(b[15]) );
  AND2X1 U94 ( .IN1(Bin[14]), .IN2(n3), .Q(b[14]) );
  AND2X1 U95 ( .IN1(Bin[13]), .IN2(n3), .Q(b[13]) );
  AND2X1 U96 ( .IN1(Bin[12]), .IN2(n3), .Q(b[12]) );
  AND2X1 U97 ( .IN1(Bin[11]), .IN2(n3), .Q(b[11]) );
  AND2X1 U98 ( .IN1(Bin[10]), .IN2(n3), .Q(b[10]) );
  AND2X1 U99 ( .IN1(Bin[0]), .IN2(n3), .Q(b[0]) );
  AND2X1 U100 ( .IN1(Ain[9]), .IN2(n3), .Q(a[9]) );
  AND2X1 U101 ( .IN1(Ain[8]), .IN2(n3), .Q(a[8]) );
  AND2X1 U102 ( .IN1(Ain[7]), .IN2(n3), .Q(a[7]) );
  AND2X1 U103 ( .IN1(Ain[6]), .IN2(n3), .Q(a[6]) );
  AND2X1 U104 ( .IN1(Ain[5]), .IN2(n3), .Q(a[5]) );
  AND2X1 U105 ( .IN1(Ain[4]), .IN2(n3), .Q(a[4]) );
  AND2X1 U106 ( .IN1(Ain[3]), .IN2(n3), .Q(a[3]) );
  AND2X1 U107 ( .IN1(Ain[2]), .IN2(n3), .Q(a[2]) );
  AND2X1 U108 ( .IN1(Ain[22]), .IN2(n3), .Q(a[22]) );
  AND2X1 U109 ( .IN1(Ain[21]), .IN2(n3), .Q(a[21]) );
  AND2X1 U110 ( .IN1(Ain[20]), .IN2(n3), .Q(a[20]) );
  AND2X1 U111 ( .IN1(Ain[1]), .IN2(n3), .Q(a[1]) );
  AND2X1 U112 ( .IN1(Ain[19]), .IN2(n3), .Q(a[19]) );
  AND2X1 U113 ( .IN1(Ain[18]), .IN2(n3), .Q(a[18]) );
  AND2X1 U114 ( .IN1(Ain[17]), .IN2(n3), .Q(a[17]) );
  AND2X1 U115 ( .IN1(Ain[16]), .IN2(n3), .Q(a[16]) );
  AND2X1 U116 ( .IN1(Ain[15]), .IN2(n3), .Q(a[15]) );
  AND2X1 U117 ( .IN1(Ain[14]), .IN2(n3), .Q(a[14]) );
  AND2X1 U118 ( .IN1(Ain[13]), .IN2(n3), .Q(a[13]) );
  AND2X1 U119 ( .IN1(Ain[12]), .IN2(n3), .Q(a[12]) );
  AND2X1 U120 ( .IN1(Ain[11]), .IN2(n3), .Q(a[11]) );
  AND2X1 U121 ( .IN1(Ain[10]), .IN2(n3), .Q(a[10]) );
  AND2X1 U122 ( .IN1(Ain[0]), .IN2(n3), .Q(a[0]) );
  MUX21X1 U123 ( .IN1(n12), .IN2(n13), .S(N24), .Q(n11) );
  AND4X1 U124 ( .IN1(n14), .IN2(N23), .IN3(N21), .IN4(N22), .Q(n13) );
  AND4X1 U125 ( .IN1(N20), .IN2(N19), .IN3(N18), .IN4(N17), .Q(n14) );
  NOR4X0 U126 ( .IN1(n15), .IN2(N17), .IN3(N19), .IN4(N18), .QN(n12) );
  OR4X1 U127 ( .IN1(N20), .IN2(N21), .IN3(N22), .IN4(N23), .Q(n15) );
  AND2X1 U128 ( .IN1(s[23]), .IN2(N69), .Q(N94) );
  MUX21X1 U129 ( .IN1(s[47]), .IN2(N68), .S(s[23]), .Q(N93) );
  MUX21X1 U130 ( .IN1(s[46]), .IN2(N67), .S(s[23]), .Q(N92) );
  MUX21X1 U131 ( .IN1(s[45]), .IN2(N66), .S(s[23]), .Q(N91) );
  MUX21X1 U132 ( .IN1(s[44]), .IN2(N65), .S(s[23]), .Q(N90) );
  MUX21X1 U133 ( .IN1(s[43]), .IN2(N64), .S(s[23]), .Q(N89) );
  MUX21X1 U134 ( .IN1(s[42]), .IN2(N63), .S(s[23]), .Q(N88) );
  MUX21X1 U135 ( .IN1(s[41]), .IN2(N62), .S(s[23]), .Q(N87) );
  MUX21X1 U136 ( .IN1(s[40]), .IN2(N61), .S(s[23]), .Q(N86) );
  MUX21X1 U137 ( .IN1(s[39]), .IN2(N60), .S(s[23]), .Q(N85) );
  MUX21X1 U138 ( .IN1(s[38]), .IN2(N59), .S(s[23]), .Q(N84) );
  MUX21X1 U139 ( .IN1(s[37]), .IN2(N58), .S(s[23]), .Q(N83) );
  MUX21X1 U140 ( .IN1(s[36]), .IN2(N57), .S(s[23]), .Q(N82) );
  MUX21X1 U141 ( .IN1(s[35]), .IN2(N56), .S(n7), .Q(N81) );
  MUX21X1 U142 ( .IN1(s[34]), .IN2(N55), .S(n7), .Q(N80) );
  MUX21X1 U143 ( .IN1(s[33]), .IN2(N54), .S(n7), .Q(N79) );
  MUX21X1 U144 ( .IN1(s[32]), .IN2(N53), .S(n7), .Q(N78) );
  MUX21X1 U145 ( .IN1(s[31]), .IN2(N52), .S(n7), .Q(N77) );
  MUX21X1 U146 ( .IN1(s[30]), .IN2(N51), .S(n7), .Q(N76) );
  MUX21X1 U147 ( .IN1(s[29]), .IN2(N50), .S(n7), .Q(N75) );
  MUX21X1 U148 ( .IN1(s[28]), .IN2(N49), .S(n7), .Q(N74) );
  MUX21X1 U149 ( .IN1(s[27]), .IN2(N48), .S(n7), .Q(N73) );
  MUX21X1 U150 ( .IN1(s[26]), .IN2(N47), .S(n7), .Q(N72) );
  MUX21X1 U151 ( .IN1(s[25]), .IN2(N46), .S(n7), .Q(N71) );
  MUX21X1 U152 ( .IN1(s[24]), .IN2(N45), .S(n7), .Q(N70) );
endmodule


module fpalu ( A, B, op, clock, reset, Result, overflow );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Result;
  input op, clock, reset;
  output overflow;
  wire   flag2, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, n1, n2, n6, net13890,
         net13888, net13894, net14211, net16090, n7, n8, n9;
  wire   [31:0] out1;
  wire   [31:0] out2;
  wire   [1:0] state;
  wire   [1:0] next_state;

  DFFARX1 \state_reg[0]  ( .D(next_state[0]), .CLK(clock), .RSTB(reset), .Q(
        state[0]), .QN(n2) );
  DFFARX1 \state_reg[1]  ( .D(next_state[1]), .CLK(clock), .RSTB(reset), .Q(
        state[1]), .QN(n1) );
  LATCHX1 \Result_reg[31]  ( .CLK(n7), .D(N53), .Q(Result[31]) );
  LATCHX1 \Result_reg[30]  ( .CLK(n7), .D(N52), .Q(Result[30]) );
  LATCHX1 \Result_reg[29]  ( .CLK(n7), .D(N51), .Q(Result[29]) );
  LATCHX1 \Result_reg[28]  ( .CLK(n7), .D(N50), .Q(Result[28]) );
  LATCHX1 \Result_reg[27]  ( .CLK(n7), .D(N49), .Q(Result[27]) );
  LATCHX1 \Result_reg[26]  ( .CLK(n7), .D(N48), .Q(Result[26]) );
  LATCHX1 \Result_reg[25]  ( .CLK(n7), .D(N47), .Q(Result[25]) );
  LATCHX1 \Result_reg[24]  ( .CLK(n7), .D(N46), .Q(Result[24]) );
  LATCHX1 \Result_reg[23]  ( .CLK(n7), .D(N45), .Q(Result[23]) );
  LATCHX1 \Result_reg[22]  ( .CLK(n7), .D(N44), .Q(Result[22]) );
  LATCHX1 \Result_reg[21]  ( .CLK(n7), .D(N43), .Q(Result[21]) );
  LATCHX1 \Result_reg[20]  ( .CLK(n7), .D(N42), .Q(Result[20]) );
  LATCHX1 \Result_reg[19]  ( .CLK(n8), .D(N41), .Q(Result[19]) );
  LATCHX1 \Result_reg[18]  ( .CLK(n8), .D(N40), .Q(Result[18]) );
  LATCHX1 \Result_reg[17]  ( .CLK(n8), .D(N39), .Q(Result[17]) );
  LATCHX1 \Result_reg[16]  ( .CLK(n8), .D(N38), .Q(Result[16]) );
  LATCHX1 \Result_reg[15]  ( .CLK(n8), .D(N37), .Q(Result[15]) );
  LATCHX1 \Result_reg[14]  ( .CLK(n8), .D(N36), .Q(Result[14]) );
  LATCHX1 \Result_reg[13]  ( .CLK(n8), .D(N35), .Q(Result[13]) );
  LATCHX1 \Result_reg[12]  ( .CLK(n8), .D(N34), .Q(Result[12]) );
  LATCHX1 \Result_reg[11]  ( .CLK(n8), .D(N33), .Q(Result[11]) );
  LATCHX1 \Result_reg[10]  ( .CLK(n8), .D(N32), .Q(Result[10]) );
  LATCHX1 \Result_reg[9]  ( .CLK(n8), .D(N31), .Q(Result[9]) );
  LATCHX1 \Result_reg[8]  ( .CLK(n8), .D(N30), .Q(Result[8]) );
  LATCHX1 \Result_reg[7]  ( .CLK(N21), .D(N29), .Q(Result[7]) );
  LATCHX1 \Result_reg[6]  ( .CLK(N21), .D(N28), .Q(Result[6]) );
  LATCHX1 \Result_reg[5]  ( .CLK(N21), .D(N27), .Q(Result[5]) );
  LATCHX1 \Result_reg[4]  ( .CLK(N21), .D(N26), .Q(Result[4]) );
  LATCHX1 \Result_reg[3]  ( .CLK(N21), .D(N25), .Q(Result[3]) );
  LATCHX1 \Result_reg[2]  ( .CLK(N21), .D(N24), .Q(Result[2]) );
  LATCHX1 \Result_reg[1]  ( .CLK(N21), .D(N23), .Q(Result[1]) );
  LATCHX1 \Result_reg[0]  ( .CLK(n8), .D(N22), .Q(Result[0]) );
  LATCHX1 overflow_reg ( .CLK(n7), .D(N54), .Q(overflow) );
  AO22X1 U10 ( .IN1(out1[31]), .IN2(net13890), .IN3(out2[31]), .IN4(net14211), 
        .Q(N53) );
  AO22X1 U11 ( .IN1(out1[30]), .IN2(net13890), .IN3(out2[30]), .IN4(n6), .Q(
        N52) );
  AO22X1 U12 ( .IN1(out1[29]), .IN2(net13890), .IN3(out2[29]), .IN4(n6), .Q(
        N51) );
  AO22X1 U13 ( .IN1(out1[28]), .IN2(net13890), .IN3(out2[28]), .IN4(net14211), 
        .Q(N50) );
  AO22X1 U14 ( .IN1(out1[27]), .IN2(net13890), .IN3(out2[27]), .IN4(net13894), 
        .Q(N49) );
  AO22X1 U15 ( .IN1(out1[26]), .IN2(net13890), .IN3(out2[26]), .IN4(net13894), 
        .Q(N48) );
  AO22X1 U16 ( .IN1(out1[25]), .IN2(net13890), .IN3(out2[25]), .IN4(net14211), 
        .Q(N47) );
  AO22X1 U17 ( .IN1(out1[24]), .IN2(net13890), .IN3(out2[24]), .IN4(n6), .Q(
        N46) );
  AO22X1 U18 ( .IN1(out1[23]), .IN2(net13890), .IN3(out2[23]), .IN4(n6), .Q(
        N45) );
  AO22X1 U19 ( .IN1(out1[22]), .IN2(net13890), .IN3(out2[22]), .IN4(net14211), 
        .Q(N44) );
  AO22X1 U20 ( .IN1(out1[21]), .IN2(net13890), .IN3(out2[21]), .IN4(net13894), 
        .Q(N43) );
  AO22X1 U21 ( .IN1(out1[20]), .IN2(net13890), .IN3(out2[20]), .IN4(net13894), 
        .Q(N42) );
  AO22X1 U22 ( .IN1(out1[19]), .IN2(net13890), .IN3(out2[19]), .IN4(net14211), 
        .Q(N41) );
  AO22X1 U23 ( .IN1(out1[18]), .IN2(net13890), .IN3(out2[18]), .IN4(n6), .Q(
        N40) );
  AO22X1 U24 ( .IN1(out1[17]), .IN2(net13888), .IN3(out2[17]), .IN4(n6), .Q(
        N39) );
  AO22X1 U25 ( .IN1(out1[16]), .IN2(net13888), .IN3(out2[16]), .IN4(net14211), 
        .Q(N38) );
  AO22X1 U26 ( .IN1(out1[15]), .IN2(net13888), .IN3(out2[15]), .IN4(net13894), 
        .Q(N37) );
  AO22X1 U27 ( .IN1(out1[14]), .IN2(net13888), .IN3(out2[14]), .IN4(net13894), 
        .Q(N36) );
  AO22X1 U28 ( .IN1(out1[13]), .IN2(net13888), .IN3(out2[13]), .IN4(net14211), 
        .Q(N35) );
  AO22X1 U29 ( .IN1(out1[12]), .IN2(net13888), .IN3(out2[12]), .IN4(n6), .Q(
        N34) );
  AO22X1 U30 ( .IN1(out1[11]), .IN2(net13888), .IN3(out2[11]), .IN4(n6), .Q(
        N33) );
  AO22X1 U31 ( .IN1(out1[10]), .IN2(net13888), .IN3(out2[10]), .IN4(net14211), 
        .Q(N32) );
  AO22X1 U32 ( .IN1(out1[9]), .IN2(net13888), .IN3(out2[9]), .IN4(net13894), 
        .Q(N31) );
  AO22X1 U33 ( .IN1(out1[8]), .IN2(net13888), .IN3(out2[8]), .IN4(net13894), 
        .Q(N30) );
  AO22X1 U34 ( .IN1(out1[7]), .IN2(net13888), .IN3(out2[7]), .IN4(net14211), 
        .Q(N29) );
  AO22X1 U35 ( .IN1(out1[6]), .IN2(net13888), .IN3(out2[6]), .IN4(n6), .Q(N28)
         );
  AO22X1 U36 ( .IN1(out1[5]), .IN2(net13888), .IN3(out2[5]), .IN4(n6), .Q(N27)
         );
  AO22X1 U37 ( .IN1(out1[4]), .IN2(net13888), .IN3(out2[4]), .IN4(net14211), 
        .Q(N26) );
  AO22X1 U38 ( .IN1(out1[3]), .IN2(net13888), .IN3(out2[3]), .IN4(net14211), 
        .Q(N25) );
  AO22X1 U39 ( .IN1(out1[2]), .IN2(net13888), .IN3(out2[2]), .IN4(net13894), 
        .Q(N24) );
  AO22X1 U40 ( .IN1(out1[1]), .IN2(net13888), .IN3(out2[1]), .IN4(n6), .Q(N23)
         );
  AO22X1 U41 ( .IN1(out1[0]), .IN2(net13888), .IN3(out2[0]), .IN4(net13894), 
        .Q(N22) );
  fpalu_add1 f1 ( .a_in(A), .b_in(B), .sum(out1) );
  fpalu_multiplier f2 ( .Ain(A), .Bin(B), .product(out2), .flag(flag2) );
  NOR2X0 U43 ( .IN1(n1), .IN2(state[0]), .QN(net13894) );
  NOR2X0 U44 ( .IN1(n1), .IN2(state[0]), .QN(net14211) );
  NAND2X1 U45 ( .IN1(state[0]), .IN2(state[1]), .QN(N21) );
  AOI21X1 U46 ( .IN1(state[1]), .IN2(state[0]), .IN3(op), .QN(next_state[0])
         );
  OA21X1 U47 ( .IN1(n1), .IN2(n2), .IN3(op), .Q(next_state[1]) );
  OR2X1 U48 ( .IN1(n2), .IN2(state[1]), .Q(net16090) );
  NOR2X0 U49 ( .IN1(n1), .IN2(state[0]), .QN(n6) );
  NBUFFX2 U50 ( .INP(N21), .Z(n8) );
  NBUFFX2 U51 ( .INP(N21), .Z(n7) );
  NAND2X1 U52 ( .IN1(net16090), .IN2(n9), .QN(N54) );
  NAND2X1 U53 ( .IN1(flag2), .IN2(net14211), .QN(n9) );
  INVX0 U54 ( .INP(net16090), .ZN(net13888) );
  INVX0 U55 ( .INP(net16090), .ZN(net13890) );
endmodule

